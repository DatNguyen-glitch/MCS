.SUBCKT dec_6to64 VDD VSS  addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] wordline[63] wordline[62] wordline[61] wordline[60] wordline[59] wordline[58] wordline[57] wordline[56] wordline[55] wordline[54] wordline[53] wordline[52] wordline[51] wordline[50] wordline[49] wordline[48] wordline[47] wordline[46] wordline[45] wordline[44] wordline[43] wordline[42] wordline[41] wordline[40] wordline[39] wordline[38] wordline[37] wordline[36] wordline[35] wordline[34] wordline[33] wordline[32] wordline[31] wordline[30] wordline[29] wordline[28] wordline[27] wordline[26] wordline[25] wordline[24] wordline[23] wordline[22] wordline[21] wordline[20] wordline[19] wordline[18] wordline[17] wordline[16] wordline[15] wordline[14] wordline[13] wordline[12] wordline[11] wordline[10] wordline[9] wordline[8] wordline[7] wordline[6] wordline[5] wordline[4] wordline[3] wordline[2] wordline[1] wordline[0]
XU88 addr[3] n33 VDD VSS  n34 NOR2xp33_ASAP7_75t_R
XU89 addr[4] VDD VSS  n23 INVx4_ASAP7_75t_R
XU90 addr[5] addr[4] VDD VSS  n33 NAND2xp5_ASAP7_75t_R
XU91 addr[5] VDD VSS  n24 INVx4_ASAP7_75t_R
XU92 addr[4] VDD VSS  n39 INVx8_ASAP7_75t_R
XU93 addr[5] VDD VSS  n36 INVx8_ASAP7_75t_R
XU94 addr[0] VDD VSS  n25 INVx8_ASAP7_75t_R
XU95 addr[2] VDD VSS  n26 INVx8_ASAP7_75t_R
XU96 addr[0] VDD VSS  n30 INVx8_ASAP7_75t_R
XU97 addr[2] VDD VSS  n29 INVx8_ASAP7_75t_R
XU98 addr[3] VDD VSS  n27 INVx8_ASAP7_75t_R
XU99 addr[3] VDD VSS  n41 INVx8_ASAP7_75t_R
XU100 addr[1] VDD VSS  n28 INVx8_ASAP7_75t_R
XU101 addr[1] VDD VSS  n31 INVx8_ASAP7_75t_R
XU102 addr[1] addr[0] addr[2] VDD VSS  n43 NOR3xp33_ASAP7_75t_R
XU103 n27 n36 n23 VDD VSS  n32 NOR3xp33_ASAP7_75t_R
XU104 n43 n32 VDD VSS  wordline[56] NAND2xp33_ASAP7_75t_R
XU105 addr[1] addr[2] n30 VDD VSS  n44 NOR3xp33_ASAP7_75t_R
XU106 n32 n44 VDD VSS  wordline[57] NAND2xp33_ASAP7_75t_R
XU107 addr[0] addr[2] n31 VDD VSS  n45 NOR3xp33_ASAP7_75t_R
XU108 n32 n45 VDD VSS  wordline[58] NAND2xp33_ASAP7_75t_R
XU109 addr[2] n25 n31 VDD VSS  n46 NOR3xp33_ASAP7_75t_R
XU110 n32 n46 VDD VSS  wordline[59] NAND2xp33_ASAP7_75t_R
XU111 addr[1] addr[0] n29 VDD VSS  n47 NOR3xp33_ASAP7_75t_R
XU112 n32 n47 VDD VSS  wordline[60] NAND2xp33_ASAP7_75t_R
XU113 addr[1] n30 n26 VDD VSS  n48 NOR3xp33_ASAP7_75t_R
XU114 n32 n48 VDD VSS  wordline[61] NAND2xp33_ASAP7_75t_R
XU115 addr[0] n28 n29 VDD VSS  n49 NOR3xp33_ASAP7_75t_R
XU116 n32 n49 VDD VSS  wordline[62] NAND2xp33_ASAP7_75t_R
XU117 n28 n25 n26 VDD VSS  n51 NOR3xp33_ASAP7_75t_R
XU118 n32 n51 VDD VSS  wordline[63] NAND2xp33_ASAP7_75t_R
XU119 n43 n34 VDD VSS  wordline[48] NAND2xp33_ASAP7_75t_R
XU120 n44 n34 VDD VSS  wordline[49] NAND2xp33_ASAP7_75t_R
XU121 n45 n34 VDD VSS  wordline[50] NAND2xp33_ASAP7_75t_R
XU122 n46 n34 VDD VSS  wordline[51] NAND2xp33_ASAP7_75t_R
XU123 n47 n34 VDD VSS  wordline[52] NAND2xp33_ASAP7_75t_R
XU124 n48 n34 VDD VSS  wordline[53] NAND2xp33_ASAP7_75t_R
XU125 n49 n34 VDD VSS  wordline[54] NAND2xp33_ASAP7_75t_R
XU126 n51 n34 VDD VSS  wordline[55] NAND2xp33_ASAP7_75t_R
XU127 addr[4] n36 n41 VDD VSS  n35 NOR3xp33_ASAP7_75t_R
XU128 n43 n35 VDD VSS  wordline[40] NAND2xp33_ASAP7_75t_R
XU129 n44 n35 VDD VSS  wordline[41] NAND2xp33_ASAP7_75t_R
XU130 n45 n35 VDD VSS  wordline[42] NAND2xp33_ASAP7_75t_R
XU131 n46 n35 VDD VSS  wordline[43] NAND2xp33_ASAP7_75t_R
XU132 n47 n35 VDD VSS  wordline[44] NAND2xp33_ASAP7_75t_R
XU133 n48 n35 VDD VSS  wordline[45] NAND2xp33_ASAP7_75t_R
XU134 n49 n35 VDD VSS  wordline[46] NAND2xp33_ASAP7_75t_R
XU135 n51 n35 VDD VSS  wordline[47] NAND2xp33_ASAP7_75t_R
XU136 addr[3] addr[4] n24 VDD VSS  n37 NOR3xp33_ASAP7_75t_R
XU137 n43 n37 VDD VSS  wordline[32] NAND2xp33_ASAP7_75t_R
XU138 n44 n37 VDD VSS  wordline[33] NAND2xp33_ASAP7_75t_R
XU139 n45 n37 VDD VSS  wordline[34] NAND2xp33_ASAP7_75t_R
XU140 n46 n37 VDD VSS  wordline[35] NAND2xp33_ASAP7_75t_R
XU141 n47 n37 VDD VSS  wordline[36] NAND2xp33_ASAP7_75t_R
XU142 n48 n37 VDD VSS  wordline[37] NAND2xp33_ASAP7_75t_R
XU143 n49 n37 VDD VSS  wordline[38] NAND2xp33_ASAP7_75t_R
XU144 n51 n37 VDD VSS  wordline[39] NAND2xp33_ASAP7_75t_R
XU145 addr[5] n27 n39 VDD VSS  n38 NOR3xp33_ASAP7_75t_R
XU146 n43 n38 VDD VSS  wordline[24] NAND2xp33_ASAP7_75t_R
XU147 n44 n38 VDD VSS  wordline[25] NAND2xp33_ASAP7_75t_R
XU148 n45 n38 VDD VSS  wordline[26] NAND2xp33_ASAP7_75t_R
XU149 n46 n38 VDD VSS  wordline[27] NAND2xp33_ASAP7_75t_R
XU150 n47 n38 VDD VSS  wordline[28] NAND2xp33_ASAP7_75t_R
XU151 n48 n38 VDD VSS  wordline[29] NAND2xp33_ASAP7_75t_R
XU152 n49 n38 VDD VSS  wordline[30] NAND2xp33_ASAP7_75t_R
XU153 n51 n38 VDD VSS  wordline[31] NAND2xp33_ASAP7_75t_R
XU154 addr[3] addr[5] n39 VDD VSS  n40 NOR3xp33_ASAP7_75t_R
XU155 n43 n40 VDD VSS  wordline[16] NAND2xp33_ASAP7_75t_R
XU156 n44 n40 VDD VSS  wordline[17] NAND2xp33_ASAP7_75t_R
XU157 n45 n40 VDD VSS  wordline[18] NAND2xp33_ASAP7_75t_R
XU158 n46 n40 VDD VSS  wordline[19] NAND2xp33_ASAP7_75t_R
XU159 n47 n40 VDD VSS  wordline[20] NAND2xp33_ASAP7_75t_R
XU160 n48 n40 VDD VSS  wordline[21] NAND2xp33_ASAP7_75t_R
XU161 n49 n40 VDD VSS  wordline[22] NAND2xp33_ASAP7_75t_R
XU162 n51 n40 VDD VSS  wordline[23] NAND2xp33_ASAP7_75t_R
XU163 addr[5] addr[4] n41 VDD VSS  n42 NOR3xp33_ASAP7_75t_R
XU164 n43 n42 VDD VSS  wordline[8] NAND2xp33_ASAP7_75t_R
XU165 n44 n42 VDD VSS  wordline[9] NAND2xp33_ASAP7_75t_R
XU166 n45 n42 VDD VSS  wordline[10] NAND2xp33_ASAP7_75t_R
XU167 n46 n42 VDD VSS  wordline[11] NAND2xp33_ASAP7_75t_R
XU168 n47 n42 VDD VSS  wordline[12] NAND2xp33_ASAP7_75t_R
XU169 n48 n42 VDD VSS  wordline[13] NAND2xp33_ASAP7_75t_R
XU170 n49 n42 VDD VSS  wordline[14] NAND2xp33_ASAP7_75t_R
XU171 n51 n42 VDD VSS  wordline[15] NAND2xp33_ASAP7_75t_R
XU172 addr[3] addr[5] addr[4] VDD VSS  n50 NOR3xp33_ASAP7_75t_R
XU173 n43 n50 VDD VSS  wordline[0] NAND2xp33_ASAP7_75t_R
XU174 n44 n50 VDD VSS  wordline[1] NAND2xp33_ASAP7_75t_R
XU175 n45 n50 VDD VSS  wordline[2] NAND2xp33_ASAP7_75t_R
XU176 n46 n50 VDD VSS  wordline[3] NAND2xp33_ASAP7_75t_R
XU177 n47 n50 VDD VSS  wordline[4] NAND2xp33_ASAP7_75t_R
XU178 n48 n50 VDD VSS  wordline[5] NAND2xp33_ASAP7_75t_R
XU179 n49 n50 VDD VSS  wordline[6] NAND2xp33_ASAP7_75t_R
XU180 n51 n50 VDD VSS  wordline[7] NAND2xp33_ASAP7_75t_R
.ENDS


