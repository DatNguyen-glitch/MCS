.SUBCKT decoder_6to64 VDD VSS  clk 
+ in_addr[5] in_addr[4] in_addr[3] in_addr[2] in_addr[1] in_addr[0] 
+ wordline[63] wordline[62] wordline[61] wordline[60] wordline[59] wordline[58] 
+ wordline[57] wordline[56] wordline[55] wordline[54] wordline[53] wordline[52] 
+ wordline[51] wordline[50] wordline[49] wordline[48] wordline[47] wordline[46] 
+ wordline[45] wordline[44] wordline[43] wordline[42] wordline[41] wordline[40] 
+ wordline[39] wordline[38] wordline[37] wordline[36] wordline[35] wordline[34] 
+ wordline[33] wordline[32] wordline[31] wordline[30] wordline[29] wordline[28] 
+ wordline[27] wordline[26] wordline[25] wordline[24] wordline[23] wordline[22] 
+ wordline[21] wordline[20] wordline[19] wordline[18] wordline[17] wordline[16] 
+ wordline[15] wordline[14] wordline[13] wordline[12] wordline[11] wordline[10] 
+ wordline[9] wordline[8] wordline[7] wordline[6] wordline[5] wordline[4] 
+ wordline[3] wordline[2] wordline[1] wordline[0]
XU90 clk VDD VSS  n46 INVx4_ASAP7_75t_SL
XU91 in_addr[0] VDD VSS  n24 INVx5_ASAP7_75t_SL
XU92 in_addr[3] VDD VSS  n25 INVx5_ASAP7_75t_SL
XU93 in_addr[4] VDD VSS  n26 INVx5_ASAP7_75t_SL
XU94 in_addr[5] VDD VSS  n27 INVx5_ASAP7_75t_SL
XU95 in_addr[1] VDD VSS  n28 INVx5_ASAP7_75t_SL
XU96 in_addr[3] VDD VSS  n29 INVx5_ASAP7_75t_SL
XU97 in_addr[3] VDD VSS  n30 INVx5_ASAP7_75t_SL
XU98 in_addr[3] VDD VSS  n39 INVx5_ASAP7_75t_SL
XU99 in_addr[0] VDD VSS  n31 INVx5_ASAP7_75t_SL
XU100 in_addr[0] VDD VSS  n32 INVx5_ASAP7_75t_SL
XU101 in_addr[4] VDD VSS  n33 INVx5_ASAP7_75t_SL
XU102 in_addr[4] VDD VSS  n34 INVx5_ASAP7_75t_SL
XU103 in_addr[0] VDD VSS  n49 INVx5_ASAP7_75t_SL
XU104 in_addr[4] VDD VSS  n40 INVx5_ASAP7_75t_SL
XU105 n61 n43 VDD VSS  wordline[6] NOR2xp67_ASAP7_75t_SL
XU106 n61 n45 VDD VSS  wordline[5] NOR2xp67_ASAP7_75t_SL
XU107 n61 n44 VDD VSS  wordline[4] NOR2xp67_ASAP7_75t_SL
XU108 n42 n51 VDD VSS  wordline[55] NOR2xp67_ASAP7_75t_SL
XU109 n42 n55 VDD VSS  wordline[47] NOR2xp67_ASAP7_75t_SL
XU110 n42 n56 VDD VSS  wordline[39] NOR2xp67_ASAP7_75t_SL
XU111 n42 n52 VDD VSS  wordline[23] NOR2xp67_ASAP7_75t_SL
XU112 n42 n53 VDD VSS  wordline[15] NOR2xp67_ASAP7_75t_SL
XU113 n42 n57 VDD VSS  wordline[31] NOR2xp67_ASAP7_75t_SL
XU114 n61 n42 VDD VSS  wordline[7] NOR2xp67_ASAP7_75t_SL
XU115 n43 n57 VDD VSS  wordline[30] NOR2xp67_ASAP7_75t_SL
XU116 n43 n53 VDD VSS  wordline[14] NOR2xp67_ASAP7_75t_SL
XU117 n43 n55 VDD VSS  wordline[46] NOR2xp67_ASAP7_75t_SL
XU118 n43 n52 VDD VSS  wordline[22] NOR2xp67_ASAP7_75t_SL
XU119 n43 n54 VDD VSS  wordline[62] NOR2xp67_ASAP7_75t_SL
XU120 n43 n56 VDD VSS  wordline[38] NOR2xp67_ASAP7_75t_SL
XU121 n44 n53 VDD VSS  wordline[12] NOR2xp67_ASAP7_75t_SL
XU122 n44 n52 VDD VSS  wordline[20] NOR2xp67_ASAP7_75t_SL
XU123 n44 n57 VDD VSS  wordline[28] NOR2xp67_ASAP7_75t_SL
XU124 n44 n51 VDD VSS  wordline[52] NOR2xp67_ASAP7_75t_SL
XU125 n44 n55 VDD VSS  wordline[44] NOR2xp67_ASAP7_75t_SL
XU126 n45 n51 VDD VSS  wordline[53] NOR2xp67_ASAP7_75t_SL
XU127 n44 n54 VDD VSS  wordline[60] NOR2xp67_ASAP7_75t_SL
XU128 n44 n56 VDD VSS  wordline[36] NOR2xp67_ASAP7_75t_SL
XU129 n45 n55 VDD VSS  wordline[45] NOR2xp67_ASAP7_75t_SL
XU130 n45 n52 VDD VSS  wordline[21] NOR2xp67_ASAP7_75t_SL
XU131 n45 n54 VDD VSS  wordline[61] NOR2xp67_ASAP7_75t_SL
XU132 n45 n57 VDD VSS  wordline[29] NOR2xp67_ASAP7_75t_SL
XU133 n45 n53 VDD VSS  wordline[13] NOR2xp67_ASAP7_75t_SL
XU134 n45 n56 VDD VSS  wordline[37] NOR2xp67_ASAP7_75t_SL
XU135 n58 n53 VDD VSS  wordline[11] NOR2xp67_ASAP7_75t_SL
XU136 n58 n52 VDD VSS  wordline[19] NOR2xp67_ASAP7_75t_SL
XU137 n58 n57 VDD VSS  wordline[27] NOR2xp67_ASAP7_75t_SL
XU138 n58 n56 VDD VSS  wordline[35] NOR2xp67_ASAP7_75t_SL
XU139 n58 n51 VDD VSS  wordline[51] NOR2xp67_ASAP7_75t_SL
XU140 n58 n54 VDD VSS  wordline[59] NOR2xp67_ASAP7_75t_SL
XU141 n47 n57 VDD VSS  wordline[24] NOR2xp67_ASAP7_75t_SL
XU142 n47 n53 VDD VSS  wordline[8] NOR2xp67_ASAP7_75t_SL
XU143 n47 n56 VDD VSS  wordline[32] NOR2xp67_ASAP7_75t_SL
XU144 n47 n52 VDD VSS  wordline[16] NOR2xp67_ASAP7_75t_SL
XU145 n47 n54 VDD VSS  wordline[56] NOR2xp67_ASAP7_75t_SL
XU146 n47 n55 VDD VSS  wordline[40] NOR2xp67_ASAP7_75t_SL
XU147 n47 n61 VDD VSS  wordline[0] NOR2xp67_ASAP7_75t_SL
XU148 n47 n51 VDD VSS  wordline[48] NOR2xp67_ASAP7_75t_SL
XU149 n59 n52 VDD VSS  wordline[17] NOR2xp67_ASAP7_75t_SL
XU150 n59 n56 VDD VSS  wordline[33] NOR2xp67_ASAP7_75t_SL
XU151 n59 n51 VDD VSS  wordline[49] NOR2xp67_ASAP7_75t_SL
XU152 n60 n51 VDD VSS  wordline[50] NOR2xp67_ASAP7_75t_SL
XU153 n59 n57 VDD VSS  wordline[25] NOR2xp67_ASAP7_75t_SL
XU154 n60 n54 VDD VSS  wordline[58] NOR2xp67_ASAP7_75t_SL
XU155 n60 n55 VDD VSS  wordline[42] NOR2xp67_ASAP7_75t_SL
XU156 n60 n52 VDD VSS  wordline[18] NOR2xp67_ASAP7_75t_SL
XU157 n60 n53 VDD VSS  wordline[10] NOR2xp67_ASAP7_75t_SL
XU158 n59 n53 VDD VSS  wordline[9] NOR2xp67_ASAP7_75t_SL
XU159 n59 n54 VDD VSS  wordline[57] NOR2xp67_ASAP7_75t_SL
XU160 n59 n55 VDD VSS  wordline[41] NOR2xp67_ASAP7_75t_SL
XU161 n60 n57 VDD VSS  wordline[26] NOR2xp67_ASAP7_75t_SL
XU162 n61 n58 VDD VSS  wordline[3] NOR2xp67_ASAP7_75t_SL
XU163 n61 n59 VDD VSS  wordline[1] NOR2xp67_ASAP7_75t_SL
XU164 n61 n60 VDD VSS  wordline[2] NOR2xp67_ASAP7_75t_SL
XU165 n42 n54 VDD VSS  wordline[63] NOR2xp67_ASAP7_75t_SL
XU166 n43 n51 VDD VSS  wordline[54] NOR2xp67_ASAP7_75t_SL
XU167 n58 n55 VDD VSS  wordline[43] NOR2xp67_ASAP7_75t_SL
XU168 n60 n56 VDD VSS  wordline[34] NOR2xp67_ASAP7_75t_SL
XU169 in_addr[5] VDD VSS  n35 INVx5_ASAP7_75t_SL
XU170 in_addr[5] VDD VSS  n36 INVx5_ASAP7_75t_SL
XU171 in_addr[5] VDD VSS  n41 INVx5_ASAP7_75t_SL
XU172 in_addr[1] VDD VSS  n37 INVx5_ASAP7_75t_SL
XU173 in_addr[1] VDD VSS  n38 INVx5_ASAP7_75t_SL
XU174 in_addr[1] VDD VSS  n48 INVx5_ASAP7_75t_SL
XU175 n35 n33 n39 VDD VSS  n61 NAND3xp33_ASAP7_75t_SL
XU176 in_addr[1] clk in_addr[2] n49 VDD VSS  n43 NAND4xp25_ASAP7_75t_SL
XU177 in_addr[0] clk in_addr[2] n48 VDD VSS  n45 NAND4xp25_ASAP7_75t_SL
XU178 clk n28 n24 in_addr[2] VDD VSS  n44 NAND4xp25_ASAP7_75t_SL
XU179 in_addr[0] in_addr[1] clk in_addr[2] VDD VSS  n42 NAND4xp25_ASAP7_75t_SL
XU180 in_addr[4] in_addr[5] n25 VDD VSS  n51 NAND3xp33_ASAP7_75t_SL
XU181 in_addr[5] in_addr[3] n26 VDD VSS  n55 NAND3xp33_ASAP7_75t_SL
XU182 in_addr[5] n34 n29 VDD VSS  n56 NAND3xp33_ASAP7_75t_SL
XU183 in_addr[5] in_addr[4] in_addr[3] VDD VSS  n54 NAND3xp33_ASAP7_75t_SL
XU184 in_addr[4] n30 n27 VDD VSS  n52 NAND3xp33_ASAP7_75t_SL
XU185 in_addr[3] n36 n40 VDD VSS  n53 NAND3xp33_ASAP7_75t_SL
XU186 in_addr[4] in_addr[3] n41 VDD VSS  n57 NAND3xp33_ASAP7_75t_SL
XU187 n46 in_addr[2] VDD VSS  n50 NOR2xp33_ASAP7_75t_SL
XU188 in_addr[0] in_addr[1] n50 VDD VSS  n58 NAND3xp33_ASAP7_75t_SL
XU189 n31 n37 n50 VDD VSS  n47 NAND3xp33_ASAP7_75t_SL
XU190 in_addr[0] n50 n38 VDD VSS  n59 NAND3xp33_ASAP7_75t_SL
XU191 in_addr[1] n50 n32 VDD VSS  n60 NAND3xp33_ASAP7_75t_SL
.ENDS


