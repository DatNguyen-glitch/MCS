.subckt sram_arr128 VDD VSS BL BLB
+ wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7]
+ wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15]
+ wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23]
+ wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31]
+ wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39]
+ wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47]
+ wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55]
+ wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63]
+ wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71]
+ wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79]
+ wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87]
+ wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95]
+ wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103]
+ wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111]
+ wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119]
+ wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
x_cell0 VDD VSS wl[0] BL BLB sram_6t
x_cell1 VDD VSS wl[1] BL BLB sram_6t
x_cell2 VDD VSS wl[2] BL BLB sram_6t
x_cell3 VDD VSS wl[3] BL BLB sram_6t
x_cell4 VDD VSS wl[4] BL BLB sram_6t
x_cell5 VDD VSS wl[5] BL BLB sram_6t
x_cell6 VDD VSS wl[6] BL BLB sram_6t
x_cell7 VDD VSS wl[7] BL BLB sram_6t
x_cell8 VDD VSS wl[8] BL BLB sram_6t
x_cell9 VDD VSS wl[9] BL BLB sram_6t
x_cell10 VDD VSS wl[10] BL BLB sram_6t
x_cell11 VDD VSS wl[11] BL BLB sram_6t
x_cell12 VDD VSS wl[12] BL BLB sram_6t
x_cell13 VDD VSS wl[13] BL BLB sram_6t
x_cell14 VDD VSS wl[14] BL BLB sram_6t
x_cell15 VDD VSS wl[15] BL BLB sram_6t
x_cell16 VDD VSS wl[16] BL BLB sram_6t
x_cell17 VDD VSS wl[17] BL BLB sram_6t
x_cell18 VDD VSS wl[18] BL BLB sram_6t
x_cell19 VDD VSS wl[19] BL BLB sram_6t
x_cell20 VDD VSS wl[20] BL BLB sram_6t
x_cell21 VDD VSS wl[21] BL BLB sram_6t
x_cell22 VDD VSS wl[22] BL BLB sram_6t
x_cell23 VDD VSS wl[23] BL BLB sram_6t
x_cell24 VDD VSS wl[24] BL BLB sram_6t
x_cell25 VDD VSS wl[25] BL BLB sram_6t
x_cell26 VDD VSS wl[26] BL BLB sram_6t
x_cell27 VDD VSS wl[27] BL BLB sram_6t
x_cell28 VDD VSS wl[28] BL BLB sram_6t
x_cell29 VDD VSS wl[29] BL BLB sram_6t
x_cell30 VDD VSS wl[30] BL BLB sram_6t
x_cell31 VDD VSS wl[31] BL BLB sram_6t
x_cell32 VDD VSS wl[32] BL BLB sram_6t
x_cell33 VDD VSS wl[33] BL BLB sram_6t
x_cell34 VDD VSS wl[34] BL BLB sram_6t
x_cell35 VDD VSS wl[35] BL BLB sram_6t
x_cell36 VDD VSS wl[36] BL BLB sram_6t
x_cell37 VDD VSS wl[37] BL BLB sram_6t
x_cell38 VDD VSS wl[38] BL BLB sram_6t
x_cell39 VDD VSS wl[39] BL BLB sram_6t
x_cell40 VDD VSS wl[40] BL BLB sram_6t
x_cell41 VDD VSS wl[41] BL BLB sram_6t
x_cell42 VDD VSS wl[42] BL BLB sram_6t
x_cell43 VDD VSS wl[43] BL BLB sram_6t
x_cell44 VDD VSS wl[44] BL BLB sram_6t
x_cell45 VDD VSS wl[45] BL BLB sram_6t
x_cell46 VDD VSS wl[46] BL BLB sram_6t
x_cell47 VDD VSS wl[47] BL BLB sram_6t
x_cell48 VDD VSS wl[48] BL BLB sram_6t
x_cell49 VDD VSS wl[49] BL BLB sram_6t
x_cell50 VDD VSS wl[50] BL BLB sram_6t
x_cell51 VDD VSS wl[51] BL BLB sram_6t
x_cell52 VDD VSS wl[52] BL BLB sram_6t
x_cell53 VDD VSS wl[53] BL BLB sram_6t
x_cell54 VDD VSS wl[54] BL BLB sram_6t
x_cell55 VDD VSS wl[55] BL BLB sram_6t
x_cell56 VDD VSS wl[56] BL BLB sram_6t
x_cell57 VDD VSS wl[57] BL BLB sram_6t
x_cell58 VDD VSS wl[58] BL BLB sram_6t
x_cell59 VDD VSS wl[59] BL BLB sram_6t
x_cell60 VDD VSS wl[60] BL BLB sram_6t
x_cell61 VDD VSS wl[61] BL BLB sram_6t
x_cell62 VDD VSS wl[62] BL BLB sram_6t
x_cell63 VDD VSS wl[63] BL BLB sram_6t
x_cell64 VDD VSS wl[64] BL BLB sram_6t
x_cell65 VDD VSS wl[65] BL BLB sram_6t
x_cell66 VDD VSS wl[66] BL BLB sram_6t
x_cell67 VDD VSS wl[67] BL BLB sram_6t
x_cell68 VDD VSS wl[68] BL BLB sram_6t
x_cell69 VDD VSS wl[69] BL BLB sram_6t
x_cell70 VDD VSS wl[70] BL BLB sram_6t
x_cell71 VDD VSS wl[71] BL BLB sram_6t
x_cell72 VDD VSS wl[72] BL BLB sram_6t
x_cell73 VDD VSS wl[73] BL BLB sram_6t
x_cell74 VDD VSS wl[74] BL BLB sram_6t
x_cell75 VDD VSS wl[75] BL BLB sram_6t
x_cell76 VDD VSS wl[76] BL BLB sram_6t
x_cell77 VDD VSS wl[77] BL BLB sram_6t
x_cell78 VDD VSS wl[78] BL BLB sram_6t
x_cell79 VDD VSS wl[79] BL BLB sram_6t
x_cell80 VDD VSS wl[80] BL BLB sram_6t
x_cell81 VDD VSS wl[81] BL BLB sram_6t
x_cell82 VDD VSS wl[82] BL BLB sram_6t
x_cell83 VDD VSS wl[83] BL BLB sram_6t
x_cell84 VDD VSS wl[84] BL BLB sram_6t
x_cell85 VDD VSS wl[85] BL BLB sram_6t
x_cell86 VDD VSS wl[86] BL BLB sram_6t
x_cell87 VDD VSS wl[87] BL BLB sram_6t
x_cell88 VDD VSS wl[88] BL BLB sram_6t
x_cell89 VDD VSS wl[89] BL BLB sram_6t
x_cell90 VDD VSS wl[90] BL BLB sram_6t
x_cell91 VDD VSS wl[91] BL BLB sram_6t
x_cell92 VDD VSS wl[92] BL BLB sram_6t
x_cell93 VDD VSS wl[93] BL BLB sram_6t
x_cell94 VDD VSS wl[94] BL BLB sram_6t
x_cell95 VDD VSS wl[95] BL BLB sram_6t
x_cell96 VDD VSS wl[96] BL BLB sram_6t
x_cell97 VDD VSS wl[97] BL BLB sram_6t
x_cell98 VDD VSS wl[98] BL BLB sram_6t
x_cell99 VDD VSS wl[99] BL BLB sram_6t
x_cell100 VDD VSS wl[100] BL BLB sram_6t
x_cell101 VDD VSS wl[101] BL BLB sram_6t
x_cell102 VDD VSS wl[102] BL BLB sram_6t
x_cell103 VDD VSS wl[103] BL BLB sram_6t
x_cell104 VDD VSS wl[104] BL BLB sram_6t
x_cell105 VDD VSS wl[105] BL BLB sram_6t
x_cell106 VDD VSS wl[106] BL BLB sram_6t
x_cell107 VDD VSS wl[107] BL BLB sram_6t
x_cell108 VDD VSS wl[108] BL BLB sram_6t
x_cell109 VDD VSS wl[109] BL BLB sram_6t
x_cell110 VDD VSS wl[110] BL BLB sram_6t
x_cell111 VDD VSS wl[111] BL BLB sram_6t
x_cell112 VDD VSS wl[112] BL BLB sram_6t
x_cell113 VDD VSS wl[113] BL BLB sram_6t
x_cell114 VDD VSS wl[114] BL BLB sram_6t
x_cell115 VDD VSS wl[115] BL BLB sram_6t
x_cell116 VDD VSS wl[116] BL BLB sram_6t
x_cell117 VDD VSS wl[117] BL BLB sram_6t
x_cell118 VDD VSS wl[118] BL BLB sram_6t
x_cell119 VDD VSS wl[119] BL BLB sram_6t
x_cell120 VDD VSS wl[120] BL BLB sram_6t
x_cell121 VDD VSS wl[121] BL BLB sram_6t
x_cell122 VDD VSS wl[122] BL BLB sram_6t
x_cell123 VDD VSS wl[123] BL BLB sram_6t
x_cell124 VDD VSS wl[124] BL BLB sram_6t
x_cell125 VDD VSS wl[125] BL BLB sram_6t
x_cell126 VDD VSS wl[126] BL BLB sram_6t
x_cell127 VDD VSS wl[127] BL BLB sram_6t
.ends
.subckt buffer_arr128 VDD VSS clk
+ in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7]
+ in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15]
+ in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23]
+ in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31]
+ in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39]
+ in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47]
+ in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55]
+ in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63]
+ in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71]
+ in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79]
+ in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87]
+ in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95]
+ in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103]
+ in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111]
+ in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119]
+ in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127]
+ out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7]
+ out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15]
+ out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23]
+ out[24] out[25] out[26] out[27] out[28] out[29] out[30] out[31]
+ out[32] out[33] out[34] out[35] out[36] out[37] out[38] out[39]
+ out[40] out[41] out[42] out[43] out[44] out[45] out[46] out[47]
+ out[48] out[49] out[50] out[51] out[52] out[53] out[54] out[55]
+ out[56] out[57] out[58] out[59] out[60] out[61] out[62] out[63]
+ out[64] out[65] out[66] out[67] out[68] out[69] out[70] out[71]
+ out[72] out[73] out[74] out[75] out[76] out[77] out[78] out[79]
+ out[80] out[81] out[82] out[83] out[84] out[85] out[86] out[87]
+ out[88] out[89] out[90] out[91] out[92] out[93] out[94] out[95]
+ out[96] out[97] out[98] out[99] out[100] out[101] out[102] out[103]
+ out[104] out[105] out[106] out[107] out[108] out[109] out[110] out[111]
+ out[112] out[113] out[114] out[115] out[116] out[117] out[118] out[119]
+ out[120] out[121] out[122] out[123] out[124] out[125] out[126] out[127]
x_buf0 VDD VSS in[0] out[0] buffer
x_and0 VSS VDD in[0] clk out[0] AND2x2_ASAP7_75t_SRAM
x_buf1 VDD VSS in[1] out[1] buffer
x_and1 VSS VDD in[1] clk out[1] AND2x2_ASAP7_75t_SRAM
x_buf2 VDD VSS in[2] out[2] buffer
x_and2 VSS VDD in[2] clk out[2] AND2x2_ASAP7_75t_SRAM
x_buf3 VDD VSS in[3] out[3] buffer
x_and3 VSS VDD in[3] clk out[3] AND2x2_ASAP7_75t_SRAM
x_buf4 VDD VSS in[4] out[4] buffer
x_and4 VSS VDD in[4] clk out[4] AND2x2_ASAP7_75t_SRAM
x_buf5 VDD VSS in[5] out[5] buffer
x_and5 VSS VDD in[5] clk out[5] AND2x2_ASAP7_75t_SRAM
x_buf6 VDD VSS in[6] out[6] buffer
x_and6 VSS VDD in[6] clk out[6] AND2x2_ASAP7_75t_SRAM
x_buf7 VDD VSS in[7] out[7] buffer
x_and7 VSS VDD in[7] clk out[7] AND2x2_ASAP7_75t_SRAM
x_buf8 VDD VSS in[8] out[8] buffer
x_and8 VSS VDD in[8] clk out[8] AND2x2_ASAP7_75t_SRAM
x_buf9 VDD VSS in[9] out[9] buffer
x_and9 VSS VDD in[9] clk out[9] AND2x2_ASAP7_75t_SRAM
x_buf10 VDD VSS in[10] out[10] buffer
x_and10 VSS VDD in[10] clk out[10] AND2x2_ASAP7_75t_SRAM
x_buf11 VDD VSS in[11] out[11] buffer
x_and11 VSS VDD in[11] clk out[11] AND2x2_ASAP7_75t_SRAM
x_buf12 VDD VSS in[12] out[12] buffer
x_and12 VSS VDD in[12] clk out[12] AND2x2_ASAP7_75t_SRAM
x_buf13 VDD VSS in[13] out[13] buffer
x_and13 VSS VDD in[13] clk out[13] AND2x2_ASAP7_75t_SRAM
x_buf14 VDD VSS in[14] out[14] buffer
x_and14 VSS VDD in[14] clk out[14] AND2x2_ASAP7_75t_SRAM
x_buf15 VDD VSS in[15] out[15] buffer
x_and15 VSS VDD in[15] clk out[15] AND2x2_ASAP7_75t_SRAM
x_buf16 VDD VSS in[16] out[16] buffer
x_and16 VSS VDD in[16] clk out[16] AND2x2_ASAP7_75t_SRAM
x_buf17 VDD VSS in[17] out[17] buffer
x_and17 VSS VDD in[17] clk out[17] AND2x2_ASAP7_75t_SRAM
x_buf18 VDD VSS in[18] out[18] buffer
x_and18 VSS VDD in[18] clk out[18] AND2x2_ASAP7_75t_SRAM
x_buf19 VDD VSS in[19] out[19] buffer
x_and19 VSS VDD in[19] clk out[19] AND2x2_ASAP7_75t_SRAM
x_buf20 VDD VSS in[20] out[20] buffer
x_and20 VSS VDD in[20] clk out[20] AND2x2_ASAP7_75t_SRAM
x_buf21 VDD VSS in[21] out[21] buffer
x_and21 VSS VDD in[21] clk out[21] AND2x2_ASAP7_75t_SRAM
x_buf22 VDD VSS in[22] out[22] buffer
x_and22 VSS VDD in[22] clk out[22] AND2x2_ASAP7_75t_SRAM
x_buf23 VDD VSS in[23] out[23] buffer
x_and23 VSS VDD in[23] clk out[23] AND2x2_ASAP7_75t_SRAM
x_buf24 VDD VSS in[24] out[24] buffer
x_and24 VSS VDD in[24] clk out[24] AND2x2_ASAP7_75t_SRAM
x_buf25 VDD VSS in[25] out[25] buffer
x_and25 VSS VDD in[25] clk out[25] AND2x2_ASAP7_75t_SRAM
x_buf26 VDD VSS in[26] out[26] buffer
x_and26 VSS VDD in[26] clk out[26] AND2x2_ASAP7_75t_SRAM
x_buf27 VDD VSS in[27] out[27] buffer
x_and27 VSS VDD in[27] clk out[27] AND2x2_ASAP7_75t_SRAM
x_buf28 VDD VSS in[28] out[28] buffer
x_and28 VSS VDD in[28] clk out[28] AND2x2_ASAP7_75t_SRAM
x_buf29 VDD VSS in[29] out[29] buffer
x_and29 VSS VDD in[29] clk out[29] AND2x2_ASAP7_75t_SRAM
x_buf30 VDD VSS in[30] out[30] buffer
x_and30 VSS VDD in[30] clk out[30] AND2x2_ASAP7_75t_SRAM
x_buf31 VDD VSS in[31] out[31] buffer
x_and31 VSS VDD in[31] clk out[31] AND2x2_ASAP7_75t_SRAM
x_buf32 VDD VSS in[32] out[32] buffer
x_and32 VSS VDD in[32] clk out[32] AND2x2_ASAP7_75t_SRAM
x_buf33 VDD VSS in[33] out[33] buffer
x_and33 VSS VDD in[33] clk out[33] AND2x2_ASAP7_75t_SRAM
x_buf34 VDD VSS in[34] out[34] buffer
x_and34 VSS VDD in[34] clk out[34] AND2x2_ASAP7_75t_SRAM
x_buf35 VDD VSS in[35] out[35] buffer
x_and35 VSS VDD in[35] clk out[35] AND2x2_ASAP7_75t_SRAM
x_buf36 VDD VSS in[36] out[36] buffer
x_and36 VSS VDD in[36] clk out[36] AND2x2_ASAP7_75t_SRAM
x_buf37 VDD VSS in[37] out[37] buffer
x_and37 VSS VDD in[37] clk out[37] AND2x2_ASAP7_75t_SRAM
x_buf38 VDD VSS in[38] out[38] buffer
x_and38 VSS VDD in[38] clk out[38] AND2x2_ASAP7_75t_SRAM
x_buf39 VDD VSS in[39] out[39] buffer
x_and39 VSS VDD in[39] clk out[39] AND2x2_ASAP7_75t_SRAM
x_buf40 VDD VSS in[40] out[40] buffer
x_and40 VSS VDD in[40] clk out[40] AND2x2_ASAP7_75t_SRAM
x_buf41 VDD VSS in[41] out[41] buffer
x_and41 VSS VDD in[41] clk out[41] AND2x2_ASAP7_75t_SRAM
x_buf42 VDD VSS in[42] out[42] buffer
x_and42 VSS VDD in[42] clk out[42] AND2x2_ASAP7_75t_SRAM
x_buf43 VDD VSS in[43] out[43] buffer
x_and43 VSS VDD in[43] clk out[43] AND2x2_ASAP7_75t_SRAM
x_buf44 VDD VSS in[44] out[44] buffer
x_and44 VSS VDD in[44] clk out[44] AND2x2_ASAP7_75t_SRAM
x_buf45 VDD VSS in[45] out[45] buffer
x_and45 VSS VDD in[45] clk out[45] AND2x2_ASAP7_75t_SRAM
x_buf46 VDD VSS in[46] out[46] buffer
x_and46 VSS VDD in[46] clk out[46] AND2x2_ASAP7_75t_SRAM
x_buf47 VDD VSS in[47] out[47] buffer
x_and47 VSS VDD in[47] clk out[47] AND2x2_ASAP7_75t_SRAM
x_buf48 VDD VSS in[48] out[48] buffer
x_and48 VSS VDD in[48] clk out[48] AND2x2_ASAP7_75t_SRAM
x_buf49 VDD VSS in[49] out[49] buffer
x_and49 VSS VDD in[49] clk out[49] AND2x2_ASAP7_75t_SRAM
x_buf50 VDD VSS in[50] out[50] buffer
x_and50 VSS VDD in[50] clk out[50] AND2x2_ASAP7_75t_SRAM
x_buf51 VDD VSS in[51] out[51] buffer
x_and51 VSS VDD in[51] clk out[51] AND2x2_ASAP7_75t_SRAM
x_buf52 VDD VSS in[52] out[52] buffer
x_and52 VSS VDD in[52] clk out[52] AND2x2_ASAP7_75t_SRAM
x_buf53 VDD VSS in[53] out[53] buffer
x_and53 VSS VDD in[53] clk out[53] AND2x2_ASAP7_75t_SRAM
x_buf54 VDD VSS in[54] out[54] buffer
x_and54 VSS VDD in[54] clk out[54] AND2x2_ASAP7_75t_SRAM
x_buf55 VDD VSS in[55] out[55] buffer
x_and55 VSS VDD in[55] clk out[55] AND2x2_ASAP7_75t_SRAM
x_buf56 VDD VSS in[56] out[56] buffer
x_and56 VSS VDD in[56] clk out[56] AND2x2_ASAP7_75t_SRAM
x_buf57 VDD VSS in[57] out[57] buffer
x_and57 VSS VDD in[57] clk out[57] AND2x2_ASAP7_75t_SRAM
x_buf58 VDD VSS in[58] out[58] buffer
x_and58 VSS VDD in[58] clk out[58] AND2x2_ASAP7_75t_SRAM
x_buf59 VDD VSS in[59] out[59] buffer
x_and59 VSS VDD in[59] clk out[59] AND2x2_ASAP7_75t_SRAM
x_buf60 VDD VSS in[60] out[60] buffer
x_and60 VSS VDD in[60] clk out[60] AND2x2_ASAP7_75t_SRAM
x_buf61 VDD VSS in[61] out[61] buffer
x_and61 VSS VDD in[61] clk out[61] AND2x2_ASAP7_75t_SRAM
x_buf62 VDD VSS in[62] out[62] buffer
x_and62 VSS VDD in[62] clk out[62] AND2x2_ASAP7_75t_SRAM
x_buf63 VDD VSS in[63] out[63] buffer
x_and63 VSS VDD in[63] clk out[63] AND2x2_ASAP7_75t_SRAM
x_buf64 VDD VSS in[64] out[64] buffer
x_and64 VSS VDD in[64] clk out[64] AND2x2_ASAP7_75t_SRAM
x_buf65 VDD VSS in[65] out[65] buffer
x_and65 VSS VDD in[65] clk out[65] AND2x2_ASAP7_75t_SRAM
x_buf66 VDD VSS in[66] out[66] buffer
x_and66 VSS VDD in[66] clk out[66] AND2x2_ASAP7_75t_SRAM
x_buf67 VDD VSS in[67] out[67] buffer
x_and67 VSS VDD in[67] clk out[67] AND2x2_ASAP7_75t_SRAM
x_buf68 VDD VSS in[68] out[68] buffer
x_and68 VSS VDD in[68] clk out[68] AND2x2_ASAP7_75t_SRAM
x_buf69 VDD VSS in[69] out[69] buffer
x_and69 VSS VDD in[69] clk out[69] AND2x2_ASAP7_75t_SRAM
x_buf70 VDD VSS in[70] out[70] buffer
x_and70 VSS VDD in[70] clk out[70] AND2x2_ASAP7_75t_SRAM
x_buf71 VDD VSS in[71] out[71] buffer
x_and71 VSS VDD in[71] clk out[71] AND2x2_ASAP7_75t_SRAM
x_buf72 VDD VSS in[72] out[72] buffer
x_and72 VSS VDD in[72] clk out[72] AND2x2_ASAP7_75t_SRAM
x_buf73 VDD VSS in[73] out[73] buffer
x_and73 VSS VDD in[73] clk out[73] AND2x2_ASAP7_75t_SRAM
x_buf74 VDD VSS in[74] out[74] buffer
x_and74 VSS VDD in[74] clk out[74] AND2x2_ASAP7_75t_SRAM
x_buf75 VDD VSS in[75] out[75] buffer
x_and75 VSS VDD in[75] clk out[75] AND2x2_ASAP7_75t_SRAM
x_buf76 VDD VSS in[76] out[76] buffer
x_and76 VSS VDD in[76] clk out[76] AND2x2_ASAP7_75t_SRAM
x_buf77 VDD VSS in[77] out[77] buffer
x_and77 VSS VDD in[77] clk out[77] AND2x2_ASAP7_75t_SRAM
x_buf78 VDD VSS in[78] out[78] buffer
x_and78 VSS VDD in[78] clk out[78] AND2x2_ASAP7_75t_SRAM
x_buf79 VDD VSS in[79] out[79] buffer
x_and79 VSS VDD in[79] clk out[79] AND2x2_ASAP7_75t_SRAM
x_buf80 VDD VSS in[80] out[80] buffer
x_and80 VSS VDD in[80] clk out[80] AND2x2_ASAP7_75t_SRAM
x_buf81 VDD VSS in[81] out[81] buffer
x_and81 VSS VDD in[81] clk out[81] AND2x2_ASAP7_75t_SRAM
x_buf82 VDD VSS in[82] out[82] buffer
x_and82 VSS VDD in[82] clk out[82] AND2x2_ASAP7_75t_SRAM
x_buf83 VDD VSS in[83] out[83] buffer
x_and83 VSS VDD in[83] clk out[83] AND2x2_ASAP7_75t_SRAM
x_buf84 VDD VSS in[84] out[84] buffer
x_and84 VSS VDD in[84] clk out[84] AND2x2_ASAP7_75t_SRAM
x_buf85 VDD VSS in[85] out[85] buffer
x_and85 VSS VDD in[85] clk out[85] AND2x2_ASAP7_75t_SRAM
x_buf86 VDD VSS in[86] out[86] buffer
x_and86 VSS VDD in[86] clk out[86] AND2x2_ASAP7_75t_SRAM
x_buf87 VDD VSS in[87] out[87] buffer
x_and87 VSS VDD in[87] clk out[87] AND2x2_ASAP7_75t_SRAM
x_buf88 VDD VSS in[88] out[88] buffer
x_and88 VSS VDD in[88] clk out[88] AND2x2_ASAP7_75t_SRAM
x_buf89 VDD VSS in[89] out[89] buffer
x_and89 VSS VDD in[89] clk out[89] AND2x2_ASAP7_75t_SRAM
x_buf90 VDD VSS in[90] out[90] buffer
x_and90 VSS VDD in[90] clk out[90] AND2x2_ASAP7_75t_SRAM
x_buf91 VDD VSS in[91] out[91] buffer
x_and91 VSS VDD in[91] clk out[91] AND2x2_ASAP7_75t_SRAM
x_buf92 VDD VSS in[92] out[92] buffer
x_and92 VSS VDD in[92] clk out[92] AND2x2_ASAP7_75t_SRAM
x_buf93 VDD VSS in[93] out[93] buffer
x_and93 VSS VDD in[93] clk out[93] AND2x2_ASAP7_75t_SRAM
x_buf94 VDD VSS in[94] out[94] buffer
x_and94 VSS VDD in[94] clk out[94] AND2x2_ASAP7_75t_SRAM
x_buf95 VDD VSS in[95] out[95] buffer
x_and95 VSS VDD in[95] clk out[95] AND2x2_ASAP7_75t_SRAM
x_buf96 VDD VSS in[96] out[96] buffer
x_and96 VSS VDD in[96] clk out[96] AND2x2_ASAP7_75t_SRAM
x_buf97 VDD VSS in[97] out[97] buffer
x_and97 VSS VDD in[97] clk out[97] AND2x2_ASAP7_75t_SRAM
x_buf98 VDD VSS in[98] out[98] buffer
x_and98 VSS VDD in[98] clk out[98] AND2x2_ASAP7_75t_SRAM
x_buf99 VDD VSS in[99] out[99] buffer
x_and99 VSS VDD in[99] clk out[99] AND2x2_ASAP7_75t_SRAM
x_buf100 VDD VSS in[100] out[100] buffer
x_and100 VSS VDD in[100] clk out[100] AND2x2_ASAP7_75t_SRAM
x_buf101 VDD VSS in[101] out[101] buffer
x_and101 VSS VDD in[101] clk out[101] AND2x2_ASAP7_75t_SRAM
x_buf102 VDD VSS in[102] out[102] buffer
x_and102 VSS VDD in[102] clk out[102] AND2x2_ASAP7_75t_SRAM
x_buf103 VDD VSS in[103] out[103] buffer
x_and103 VSS VDD in[103] clk out[103] AND2x2_ASAP7_75t_SRAM
x_buf104 VDD VSS in[104] out[104] buffer
x_and104 VSS VDD in[104] clk out[104] AND2x2_ASAP7_75t_SRAM
x_buf105 VDD VSS in[105] out[105] buffer
x_and105 VSS VDD in[105] clk out[105] AND2x2_ASAP7_75t_SRAM
x_buf106 VDD VSS in[106] out[106] buffer
x_and106 VSS VDD in[106] clk out[106] AND2x2_ASAP7_75t_SRAM
x_buf107 VDD VSS in[107] out[107] buffer
x_and107 VSS VDD in[107] clk out[107] AND2x2_ASAP7_75t_SRAM
x_buf108 VDD VSS in[108] out[108] buffer
x_and108 VSS VDD in[108] clk out[108] AND2x2_ASAP7_75t_SRAM
x_buf109 VDD VSS in[109] out[109] buffer
x_and109 VSS VDD in[109] clk out[109] AND2x2_ASAP7_75t_SRAM
x_buf110 VDD VSS in[110] out[110] buffer
x_and110 VSS VDD in[110] clk out[110] AND2x2_ASAP7_75t_SRAM
x_buf111 VDD VSS in[111] out[111] buffer
x_and111 VSS VDD in[111] clk out[111] AND2x2_ASAP7_75t_SRAM
x_buf112 VDD VSS in[112] out[112] buffer
x_and112 VSS VDD in[112] clk out[112] AND2x2_ASAP7_75t_SRAM
x_buf113 VDD VSS in[113] out[113] buffer
x_and113 VSS VDD in[113] clk out[113] AND2x2_ASAP7_75t_SRAM
x_buf114 VDD VSS in[114] out[114] buffer
x_and114 VSS VDD in[114] clk out[114] AND2x2_ASAP7_75t_SRAM
x_buf115 VDD VSS in[115] out[115] buffer
x_and115 VSS VDD in[115] clk out[115] AND2x2_ASAP7_75t_SRAM
x_buf116 VDD VSS in[116] out[116] buffer
x_and116 VSS VDD in[116] clk out[116] AND2x2_ASAP7_75t_SRAM
x_buf117 VDD VSS in[117] out[117] buffer
x_and117 VSS VDD in[117] clk out[117] AND2x2_ASAP7_75t_SRAM
x_buf118 VDD VSS in[118] out[118] buffer
x_and118 VSS VDD in[118] clk out[118] AND2x2_ASAP7_75t_SRAM
x_buf119 VDD VSS in[119] out[119] buffer
x_and119 VSS VDD in[119] clk out[119] AND2x2_ASAP7_75t_SRAM
x_buf120 VDD VSS in[120] out[120] buffer
x_and120 VSS VDD in[120] clk out[120] AND2x2_ASAP7_75t_SRAM
x_buf121 VDD VSS in[121] out[121] buffer
x_and121 VSS VDD in[121] clk out[121] AND2x2_ASAP7_75t_SRAM
x_buf122 VDD VSS in[122] out[122] buffer
x_and122 VSS VDD in[122] clk out[122] AND2x2_ASAP7_75t_SRAM
x_buf123 VDD VSS in[123] out[123] buffer
x_and123 VSS VDD in[123] clk out[123] AND2x2_ASAP7_75t_SRAM
x_buf124 VDD VSS in[124] out[124] buffer
x_and124 VSS VDD in[124] clk out[124] AND2x2_ASAP7_75t_SRAM
x_buf125 VDD VSS in[125] out[125] buffer
x_and125 VSS VDD in[125] clk out[125] AND2x2_ASAP7_75t_SRAM
x_buf126 VDD VSS in[126] out[126] buffer
x_and126 VSS VDD in[126] clk out[126] AND2x2_ASAP7_75t_SRAM
x_buf127 VDD VSS in[127] out[127] buffer
x_and127 VSS VDD in[127] clk out[127] AND2x2_ASAP7_75t_SRAM
.ends
.nodeset v(x_sram_arr0.x_cell0.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell1.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell2.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell3.q) = 0
.nodeset v(x_sram_arr0.x_cell4.q) = 0
.nodeset v(x_sram_arr0.x_cell5.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell6.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell7.q) = 0
.nodeset v(x_sram_arr0.x_cell8.q) = 0
.nodeset v(x_sram_arr0.x_cell9.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell10.q) = 0
.nodeset v(x_sram_arr0.x_cell11.q) = 0
.nodeset v(x_sram_arr0.x_cell12.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell13.q) = 0
.nodeset v(x_sram_arr0.x_cell14.q) = 0
.nodeset v(x_sram_arr0.x_cell15.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell16.q) = 0
.nodeset v(x_sram_arr0.x_cell17.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell18.q) = 0
.nodeset v(x_sram_arr0.x_cell19.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell20.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell21.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell22.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell23.q) = 0
.nodeset v(x_sram_arr0.x_cell24.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell25.q) = 0
.nodeset v(x_sram_arr0.x_cell26.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell27.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell28.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell29.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell30.q) = 0
.nodeset v(x_sram_arr0.x_cell31.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell32.q) = 0
.nodeset v(x_sram_arr0.x_cell33.q) = 0
.nodeset v(x_sram_arr0.x_cell34.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell35.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell36.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell37.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell38.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell39.q) = 0
.nodeset v(x_sram_arr0.x_cell40.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell41.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell42.q) = 0
.nodeset v(x_sram_arr0.x_cell43.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell44.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell45.q) = 0
.nodeset v(x_sram_arr0.x_cell46.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell47.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell48.q) = 0
.nodeset v(x_sram_arr0.x_cell49.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell50.q) = 0
.nodeset v(x_sram_arr0.x_cell51.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell52.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell53.q) = 0
.nodeset v(x_sram_arr0.x_cell54.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell55.q) = 0
.nodeset v(x_sram_arr0.x_cell56.q) = 0
.nodeset v(x_sram_arr0.x_cell57.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell58.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell59.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell60.q) = 0
.nodeset v(x_sram_arr0.x_cell61.q) = 0
.nodeset v(x_sram_arr0.x_cell62.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell63.q) = 0
.nodeset v(x_sram_arr0.x_cell64.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell65.q) = 0
.nodeset v(x_sram_arr0.x_cell66.q) = 0
.nodeset v(x_sram_arr0.x_cell67.q) = 0
.nodeset v(x_sram_arr0.x_cell68.q) = 0
.nodeset v(x_sram_arr0.x_cell69.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell70.q) = 0
.nodeset v(x_sram_arr0.x_cell71.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell72.q) = 0
.nodeset v(x_sram_arr0.x_cell73.q) = 0
.nodeset v(x_sram_arr0.x_cell74.q) = 0
.nodeset v(x_sram_arr0.x_cell75.q) = 0
.nodeset v(x_sram_arr0.x_cell76.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell77.q) = 0
.nodeset v(x_sram_arr0.x_cell78.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell79.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell80.q) = 0
.nodeset v(x_sram_arr0.x_cell81.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell82.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell83.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell84.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell85.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell86.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell87.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell88.q) = 0
.nodeset v(x_sram_arr0.x_cell89.q) = 0
.nodeset v(x_sram_arr0.x_cell90.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell91.q) = 0
.nodeset v(x_sram_arr0.x_cell92.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell93.q) = 0
.nodeset v(x_sram_arr0.x_cell94.q) = 0
.nodeset v(x_sram_arr0.x_cell95.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell96.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell97.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell98.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell99.q) = 0
.nodeset v(x_sram_arr0.x_cell100.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell101.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell102.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell103.q) = 0
.nodeset v(x_sram_arr0.x_cell104.q) = 0
.nodeset v(x_sram_arr0.x_cell105.q) = 0
.nodeset v(x_sram_arr0.x_cell106.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell107.q) = 0
.nodeset v(x_sram_arr0.x_cell108.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell109.q) = 0
.nodeset v(x_sram_arr0.x_cell110.q) = 0
.nodeset v(x_sram_arr0.x_cell111.q) = 0
.nodeset v(x_sram_arr0.x_cell112.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell113.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell114.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell115.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell116.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell117.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell118.q) = 0
.nodeset v(x_sram_arr0.x_cell119.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell120.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell121.q) = 0
.nodeset v(x_sram_arr0.x_cell122.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell123.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell124.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell125.q) = 0
.nodeset v(x_sram_arr0.x_cell126.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell127.q) = 0
