.subckt sram_arr512 VDD VSS BL BLB
+ wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7]
+ wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15]
+ wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23]
+ wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31]
+ wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39]
+ wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47]
+ wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55]
+ wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63]
+ wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71]
+ wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79]
+ wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87]
+ wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95]
+ wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103]
+ wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111]
+ wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119]
+ wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
+ wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135]
+ wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143]
+ wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151]
+ wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159]
+ wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167]
+ wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175]
+ wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183]
+ wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191]
+ wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199]
+ wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207]
+ wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215]
+ wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223]
+ wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231]
+ wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239]
+ wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247]
+ wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255]
+ wl[256] wl[257] wl[258] wl[259] wl[260] wl[261] wl[262] wl[263]
+ wl[264] wl[265] wl[266] wl[267] wl[268] wl[269] wl[270] wl[271]
+ wl[272] wl[273] wl[274] wl[275] wl[276] wl[277] wl[278] wl[279]
+ wl[280] wl[281] wl[282] wl[283] wl[284] wl[285] wl[286] wl[287]
+ wl[288] wl[289] wl[290] wl[291] wl[292] wl[293] wl[294] wl[295]
+ wl[296] wl[297] wl[298] wl[299] wl[300] wl[301] wl[302] wl[303]
+ wl[304] wl[305] wl[306] wl[307] wl[308] wl[309] wl[310] wl[311]
+ wl[312] wl[313] wl[314] wl[315] wl[316] wl[317] wl[318] wl[319]
+ wl[320] wl[321] wl[322] wl[323] wl[324] wl[325] wl[326] wl[327]
+ wl[328] wl[329] wl[330] wl[331] wl[332] wl[333] wl[334] wl[335]
+ wl[336] wl[337] wl[338] wl[339] wl[340] wl[341] wl[342] wl[343]
+ wl[344] wl[345] wl[346] wl[347] wl[348] wl[349] wl[350] wl[351]
+ wl[352] wl[353] wl[354] wl[355] wl[356] wl[357] wl[358] wl[359]
+ wl[360] wl[361] wl[362] wl[363] wl[364] wl[365] wl[366] wl[367]
+ wl[368] wl[369] wl[370] wl[371] wl[372] wl[373] wl[374] wl[375]
+ wl[376] wl[377] wl[378] wl[379] wl[380] wl[381] wl[382] wl[383]
+ wl[384] wl[385] wl[386] wl[387] wl[388] wl[389] wl[390] wl[391]
+ wl[392] wl[393] wl[394] wl[395] wl[396] wl[397] wl[398] wl[399]
+ wl[400] wl[401] wl[402] wl[403] wl[404] wl[405] wl[406] wl[407]
+ wl[408] wl[409] wl[410] wl[411] wl[412] wl[413] wl[414] wl[415]
+ wl[416] wl[417] wl[418] wl[419] wl[420] wl[421] wl[422] wl[423]
+ wl[424] wl[425] wl[426] wl[427] wl[428] wl[429] wl[430] wl[431]
+ wl[432] wl[433] wl[434] wl[435] wl[436] wl[437] wl[438] wl[439]
+ wl[440] wl[441] wl[442] wl[443] wl[444] wl[445] wl[446] wl[447]
+ wl[448] wl[449] wl[450] wl[451] wl[452] wl[453] wl[454] wl[455]
+ wl[456] wl[457] wl[458] wl[459] wl[460] wl[461] wl[462] wl[463]
+ wl[464] wl[465] wl[466] wl[467] wl[468] wl[469] wl[470] wl[471]
+ wl[472] wl[473] wl[474] wl[475] wl[476] wl[477] wl[478] wl[479]
+ wl[480] wl[481] wl[482] wl[483] wl[484] wl[485] wl[486] wl[487]
+ wl[488] wl[489] wl[490] wl[491] wl[492] wl[493] wl[494] wl[495]
+ wl[496] wl[497] wl[498] wl[499] wl[500] wl[501] wl[502] wl[503]
+ wl[504] wl[505] wl[506] wl[507] wl[508] wl[509] wl[510] wl[511]
x_cell0 VDD VSS wl[0] BL BLB sram_6t
x_cell1 VDD VSS wl[1] BL BLB sram_6t
x_cell2 VDD VSS wl[2] BL BLB sram_6t
x_cell3 VDD VSS wl[3] BL BLB sram_6t
x_cell4 VDD VSS wl[4] BL BLB sram_6t
x_cell5 VDD VSS wl[5] BL BLB sram_6t
x_cell6 VDD VSS wl[6] BL BLB sram_6t
x_cell7 VDD VSS wl[7] BL BLB sram_6t
x_cell8 VDD VSS wl[8] BL BLB sram_6t
x_cell9 VDD VSS wl[9] BL BLB sram_6t
x_cell10 VDD VSS wl[10] BL BLB sram_6t
x_cell11 VDD VSS wl[11] BL BLB sram_6t
x_cell12 VDD VSS wl[12] BL BLB sram_6t
x_cell13 VDD VSS wl[13] BL BLB sram_6t
x_cell14 VDD VSS wl[14] BL BLB sram_6t
x_cell15 VDD VSS wl[15] BL BLB sram_6t
x_cell16 VDD VSS wl[16] BL BLB sram_6t
x_cell17 VDD VSS wl[17] BL BLB sram_6t
x_cell18 VDD VSS wl[18] BL BLB sram_6t
x_cell19 VDD VSS wl[19] BL BLB sram_6t
x_cell20 VDD VSS wl[20] BL BLB sram_6t
x_cell21 VDD VSS wl[21] BL BLB sram_6t
x_cell22 VDD VSS wl[22] BL BLB sram_6t
x_cell23 VDD VSS wl[23] BL BLB sram_6t
x_cell24 VDD VSS wl[24] BL BLB sram_6t
x_cell25 VDD VSS wl[25] BL BLB sram_6t
x_cell26 VDD VSS wl[26] BL BLB sram_6t
x_cell27 VDD VSS wl[27] BL BLB sram_6t
x_cell28 VDD VSS wl[28] BL BLB sram_6t
x_cell29 VDD VSS wl[29] BL BLB sram_6t
x_cell30 VDD VSS wl[30] BL BLB sram_6t
x_cell31 VDD VSS wl[31] BL BLB sram_6t
x_cell32 VDD VSS wl[32] BL BLB sram_6t
x_cell33 VDD VSS wl[33] BL BLB sram_6t
x_cell34 VDD VSS wl[34] BL BLB sram_6t
x_cell35 VDD VSS wl[35] BL BLB sram_6t
x_cell36 VDD VSS wl[36] BL BLB sram_6t
x_cell37 VDD VSS wl[37] BL BLB sram_6t
x_cell38 VDD VSS wl[38] BL BLB sram_6t
x_cell39 VDD VSS wl[39] BL BLB sram_6t
x_cell40 VDD VSS wl[40] BL BLB sram_6t
x_cell41 VDD VSS wl[41] BL BLB sram_6t
x_cell42 VDD VSS wl[42] BL BLB sram_6t
x_cell43 VDD VSS wl[43] BL BLB sram_6t
x_cell44 VDD VSS wl[44] BL BLB sram_6t
x_cell45 VDD VSS wl[45] BL BLB sram_6t
x_cell46 VDD VSS wl[46] BL BLB sram_6t
x_cell47 VDD VSS wl[47] BL BLB sram_6t
x_cell48 VDD VSS wl[48] BL BLB sram_6t
x_cell49 VDD VSS wl[49] BL BLB sram_6t
x_cell50 VDD VSS wl[50] BL BLB sram_6t
x_cell51 VDD VSS wl[51] BL BLB sram_6t
x_cell52 VDD VSS wl[52] BL BLB sram_6t
x_cell53 VDD VSS wl[53] BL BLB sram_6t
x_cell54 VDD VSS wl[54] BL BLB sram_6t
x_cell55 VDD VSS wl[55] BL BLB sram_6t
x_cell56 VDD VSS wl[56] BL BLB sram_6t
x_cell57 VDD VSS wl[57] BL BLB sram_6t
x_cell58 VDD VSS wl[58] BL BLB sram_6t
x_cell59 VDD VSS wl[59] BL BLB sram_6t
x_cell60 VDD VSS wl[60] BL BLB sram_6t
x_cell61 VDD VSS wl[61] BL BLB sram_6t
x_cell62 VDD VSS wl[62] BL BLB sram_6t
x_cell63 VDD VSS wl[63] BL BLB sram_6t
x_cell64 VDD VSS wl[64] BL BLB sram_6t
x_cell65 VDD VSS wl[65] BL BLB sram_6t
x_cell66 VDD VSS wl[66] BL BLB sram_6t
x_cell67 VDD VSS wl[67] BL BLB sram_6t
x_cell68 VDD VSS wl[68] BL BLB sram_6t
x_cell69 VDD VSS wl[69] BL BLB sram_6t
x_cell70 VDD VSS wl[70] BL BLB sram_6t
x_cell71 VDD VSS wl[71] BL BLB sram_6t
x_cell72 VDD VSS wl[72] BL BLB sram_6t
x_cell73 VDD VSS wl[73] BL BLB sram_6t
x_cell74 VDD VSS wl[74] BL BLB sram_6t
x_cell75 VDD VSS wl[75] BL BLB sram_6t
x_cell76 VDD VSS wl[76] BL BLB sram_6t
x_cell77 VDD VSS wl[77] BL BLB sram_6t
x_cell78 VDD VSS wl[78] BL BLB sram_6t
x_cell79 VDD VSS wl[79] BL BLB sram_6t
x_cell80 VDD VSS wl[80] BL BLB sram_6t
x_cell81 VDD VSS wl[81] BL BLB sram_6t
x_cell82 VDD VSS wl[82] BL BLB sram_6t
x_cell83 VDD VSS wl[83] BL BLB sram_6t
x_cell84 VDD VSS wl[84] BL BLB sram_6t
x_cell85 VDD VSS wl[85] BL BLB sram_6t
x_cell86 VDD VSS wl[86] BL BLB sram_6t
x_cell87 VDD VSS wl[87] BL BLB sram_6t
x_cell88 VDD VSS wl[88] BL BLB sram_6t
x_cell89 VDD VSS wl[89] BL BLB sram_6t
x_cell90 VDD VSS wl[90] BL BLB sram_6t
x_cell91 VDD VSS wl[91] BL BLB sram_6t
x_cell92 VDD VSS wl[92] BL BLB sram_6t
x_cell93 VDD VSS wl[93] BL BLB sram_6t
x_cell94 VDD VSS wl[94] BL BLB sram_6t
x_cell95 VDD VSS wl[95] BL BLB sram_6t
x_cell96 VDD VSS wl[96] BL BLB sram_6t
x_cell97 VDD VSS wl[97] BL BLB sram_6t
x_cell98 VDD VSS wl[98] BL BLB sram_6t
x_cell99 VDD VSS wl[99] BL BLB sram_6t
x_cell100 VDD VSS wl[100] BL BLB sram_6t
x_cell101 VDD VSS wl[101] BL BLB sram_6t
x_cell102 VDD VSS wl[102] BL BLB sram_6t
x_cell103 VDD VSS wl[103] BL BLB sram_6t
x_cell104 VDD VSS wl[104] BL BLB sram_6t
x_cell105 VDD VSS wl[105] BL BLB sram_6t
x_cell106 VDD VSS wl[106] BL BLB sram_6t
x_cell107 VDD VSS wl[107] BL BLB sram_6t
x_cell108 VDD VSS wl[108] BL BLB sram_6t
x_cell109 VDD VSS wl[109] BL BLB sram_6t
x_cell110 VDD VSS wl[110] BL BLB sram_6t
x_cell111 VDD VSS wl[111] BL BLB sram_6t
x_cell112 VDD VSS wl[112] BL BLB sram_6t
x_cell113 VDD VSS wl[113] BL BLB sram_6t
x_cell114 VDD VSS wl[114] BL BLB sram_6t
x_cell115 VDD VSS wl[115] BL BLB sram_6t
x_cell116 VDD VSS wl[116] BL BLB sram_6t
x_cell117 VDD VSS wl[117] BL BLB sram_6t
x_cell118 VDD VSS wl[118] BL BLB sram_6t
x_cell119 VDD VSS wl[119] BL BLB sram_6t
x_cell120 VDD VSS wl[120] BL BLB sram_6t
x_cell121 VDD VSS wl[121] BL BLB sram_6t
x_cell122 VDD VSS wl[122] BL BLB sram_6t
x_cell123 VDD VSS wl[123] BL BLB sram_6t
x_cell124 VDD VSS wl[124] BL BLB sram_6t
x_cell125 VDD VSS wl[125] BL BLB sram_6t
x_cell126 VDD VSS wl[126] BL BLB sram_6t
x_cell127 VDD VSS wl[127] BL BLB sram_6t
x_cell128 VDD VSS wl[128] BL BLB sram_6t
x_cell129 VDD VSS wl[129] BL BLB sram_6t
x_cell130 VDD VSS wl[130] BL BLB sram_6t
x_cell131 VDD VSS wl[131] BL BLB sram_6t
x_cell132 VDD VSS wl[132] BL BLB sram_6t
x_cell133 VDD VSS wl[133] BL BLB sram_6t
x_cell134 VDD VSS wl[134] BL BLB sram_6t
x_cell135 VDD VSS wl[135] BL BLB sram_6t
x_cell136 VDD VSS wl[136] BL BLB sram_6t
x_cell137 VDD VSS wl[137] BL BLB sram_6t
x_cell138 VDD VSS wl[138] BL BLB sram_6t
x_cell139 VDD VSS wl[139] BL BLB sram_6t
x_cell140 VDD VSS wl[140] BL BLB sram_6t
x_cell141 VDD VSS wl[141] BL BLB sram_6t
x_cell142 VDD VSS wl[142] BL BLB sram_6t
x_cell143 VDD VSS wl[143] BL BLB sram_6t
x_cell144 VDD VSS wl[144] BL BLB sram_6t
x_cell145 VDD VSS wl[145] BL BLB sram_6t
x_cell146 VDD VSS wl[146] BL BLB sram_6t
x_cell147 VDD VSS wl[147] BL BLB sram_6t
x_cell148 VDD VSS wl[148] BL BLB sram_6t
x_cell149 VDD VSS wl[149] BL BLB sram_6t
x_cell150 VDD VSS wl[150] BL BLB sram_6t
x_cell151 VDD VSS wl[151] BL BLB sram_6t
x_cell152 VDD VSS wl[152] BL BLB sram_6t
x_cell153 VDD VSS wl[153] BL BLB sram_6t
x_cell154 VDD VSS wl[154] BL BLB sram_6t
x_cell155 VDD VSS wl[155] BL BLB sram_6t
x_cell156 VDD VSS wl[156] BL BLB sram_6t
x_cell157 VDD VSS wl[157] BL BLB sram_6t
x_cell158 VDD VSS wl[158] BL BLB sram_6t
x_cell159 VDD VSS wl[159] BL BLB sram_6t
x_cell160 VDD VSS wl[160] BL BLB sram_6t
x_cell161 VDD VSS wl[161] BL BLB sram_6t
x_cell162 VDD VSS wl[162] BL BLB sram_6t
x_cell163 VDD VSS wl[163] BL BLB sram_6t
x_cell164 VDD VSS wl[164] BL BLB sram_6t
x_cell165 VDD VSS wl[165] BL BLB sram_6t
x_cell166 VDD VSS wl[166] BL BLB sram_6t
x_cell167 VDD VSS wl[167] BL BLB sram_6t
x_cell168 VDD VSS wl[168] BL BLB sram_6t
x_cell169 VDD VSS wl[169] BL BLB sram_6t
x_cell170 VDD VSS wl[170] BL BLB sram_6t
x_cell171 VDD VSS wl[171] BL BLB sram_6t
x_cell172 VDD VSS wl[172] BL BLB sram_6t
x_cell173 VDD VSS wl[173] BL BLB sram_6t
x_cell174 VDD VSS wl[174] BL BLB sram_6t
x_cell175 VDD VSS wl[175] BL BLB sram_6t
x_cell176 VDD VSS wl[176] BL BLB sram_6t
x_cell177 VDD VSS wl[177] BL BLB sram_6t
x_cell178 VDD VSS wl[178] BL BLB sram_6t
x_cell179 VDD VSS wl[179] BL BLB sram_6t
x_cell180 VDD VSS wl[180] BL BLB sram_6t
x_cell181 VDD VSS wl[181] BL BLB sram_6t
x_cell182 VDD VSS wl[182] BL BLB sram_6t
x_cell183 VDD VSS wl[183] BL BLB sram_6t
x_cell184 VDD VSS wl[184] BL BLB sram_6t
x_cell185 VDD VSS wl[185] BL BLB sram_6t
x_cell186 VDD VSS wl[186] BL BLB sram_6t
x_cell187 VDD VSS wl[187] BL BLB sram_6t
x_cell188 VDD VSS wl[188] BL BLB sram_6t
x_cell189 VDD VSS wl[189] BL BLB sram_6t
x_cell190 VDD VSS wl[190] BL BLB sram_6t
x_cell191 VDD VSS wl[191] BL BLB sram_6t
x_cell192 VDD VSS wl[192] BL BLB sram_6t
x_cell193 VDD VSS wl[193] BL BLB sram_6t
x_cell194 VDD VSS wl[194] BL BLB sram_6t
x_cell195 VDD VSS wl[195] BL BLB sram_6t
x_cell196 VDD VSS wl[196] BL BLB sram_6t
x_cell197 VDD VSS wl[197] BL BLB sram_6t
x_cell198 VDD VSS wl[198] BL BLB sram_6t
x_cell199 VDD VSS wl[199] BL BLB sram_6t
x_cell200 VDD VSS wl[200] BL BLB sram_6t
x_cell201 VDD VSS wl[201] BL BLB sram_6t
x_cell202 VDD VSS wl[202] BL BLB sram_6t
x_cell203 VDD VSS wl[203] BL BLB sram_6t
x_cell204 VDD VSS wl[204] BL BLB sram_6t
x_cell205 VDD VSS wl[205] BL BLB sram_6t
x_cell206 VDD VSS wl[206] BL BLB sram_6t
x_cell207 VDD VSS wl[207] BL BLB sram_6t
x_cell208 VDD VSS wl[208] BL BLB sram_6t
x_cell209 VDD VSS wl[209] BL BLB sram_6t
x_cell210 VDD VSS wl[210] BL BLB sram_6t
x_cell211 VDD VSS wl[211] BL BLB sram_6t
x_cell212 VDD VSS wl[212] BL BLB sram_6t
x_cell213 VDD VSS wl[213] BL BLB sram_6t
x_cell214 VDD VSS wl[214] BL BLB sram_6t
x_cell215 VDD VSS wl[215] BL BLB sram_6t
x_cell216 VDD VSS wl[216] BL BLB sram_6t
x_cell217 VDD VSS wl[217] BL BLB sram_6t
x_cell218 VDD VSS wl[218] BL BLB sram_6t
x_cell219 VDD VSS wl[219] BL BLB sram_6t
x_cell220 VDD VSS wl[220] BL BLB sram_6t
x_cell221 VDD VSS wl[221] BL BLB sram_6t
x_cell222 VDD VSS wl[222] BL BLB sram_6t
x_cell223 VDD VSS wl[223] BL BLB sram_6t
x_cell224 VDD VSS wl[224] BL BLB sram_6t
x_cell225 VDD VSS wl[225] BL BLB sram_6t
x_cell226 VDD VSS wl[226] BL BLB sram_6t
x_cell227 VDD VSS wl[227] BL BLB sram_6t
x_cell228 VDD VSS wl[228] BL BLB sram_6t
x_cell229 VDD VSS wl[229] BL BLB sram_6t
x_cell230 VDD VSS wl[230] BL BLB sram_6t
x_cell231 VDD VSS wl[231] BL BLB sram_6t
x_cell232 VDD VSS wl[232] BL BLB sram_6t
x_cell233 VDD VSS wl[233] BL BLB sram_6t
x_cell234 VDD VSS wl[234] BL BLB sram_6t
x_cell235 VDD VSS wl[235] BL BLB sram_6t
x_cell236 VDD VSS wl[236] BL BLB sram_6t
x_cell237 VDD VSS wl[237] BL BLB sram_6t
x_cell238 VDD VSS wl[238] BL BLB sram_6t
x_cell239 VDD VSS wl[239] BL BLB sram_6t
x_cell240 VDD VSS wl[240] BL BLB sram_6t
x_cell241 VDD VSS wl[241] BL BLB sram_6t
x_cell242 VDD VSS wl[242] BL BLB sram_6t
x_cell243 VDD VSS wl[243] BL BLB sram_6t
x_cell244 VDD VSS wl[244] BL BLB sram_6t
x_cell245 VDD VSS wl[245] BL BLB sram_6t
x_cell246 VDD VSS wl[246] BL BLB sram_6t
x_cell247 VDD VSS wl[247] BL BLB sram_6t
x_cell248 VDD VSS wl[248] BL BLB sram_6t
x_cell249 VDD VSS wl[249] BL BLB sram_6t
x_cell250 VDD VSS wl[250] BL BLB sram_6t
x_cell251 VDD VSS wl[251] BL BLB sram_6t
x_cell252 VDD VSS wl[252] BL BLB sram_6t
x_cell253 VDD VSS wl[253] BL BLB sram_6t
x_cell254 VDD VSS wl[254] BL BLB sram_6t
x_cell255 VDD VSS wl[255] BL BLB sram_6t
x_cell256 VDD VSS wl[256] BL BLB sram_6t
x_cell257 VDD VSS wl[257] BL BLB sram_6t
x_cell258 VDD VSS wl[258] BL BLB sram_6t
x_cell259 VDD VSS wl[259] BL BLB sram_6t
x_cell260 VDD VSS wl[260] BL BLB sram_6t
x_cell261 VDD VSS wl[261] BL BLB sram_6t
x_cell262 VDD VSS wl[262] BL BLB sram_6t
x_cell263 VDD VSS wl[263] BL BLB sram_6t
x_cell264 VDD VSS wl[264] BL BLB sram_6t
x_cell265 VDD VSS wl[265] BL BLB sram_6t
x_cell266 VDD VSS wl[266] BL BLB sram_6t
x_cell267 VDD VSS wl[267] BL BLB sram_6t
x_cell268 VDD VSS wl[268] BL BLB sram_6t
x_cell269 VDD VSS wl[269] BL BLB sram_6t
x_cell270 VDD VSS wl[270] BL BLB sram_6t
x_cell271 VDD VSS wl[271] BL BLB sram_6t
x_cell272 VDD VSS wl[272] BL BLB sram_6t
x_cell273 VDD VSS wl[273] BL BLB sram_6t
x_cell274 VDD VSS wl[274] BL BLB sram_6t
x_cell275 VDD VSS wl[275] BL BLB sram_6t
x_cell276 VDD VSS wl[276] BL BLB sram_6t
x_cell277 VDD VSS wl[277] BL BLB sram_6t
x_cell278 VDD VSS wl[278] BL BLB sram_6t
x_cell279 VDD VSS wl[279] BL BLB sram_6t
x_cell280 VDD VSS wl[280] BL BLB sram_6t
x_cell281 VDD VSS wl[281] BL BLB sram_6t
x_cell282 VDD VSS wl[282] BL BLB sram_6t
x_cell283 VDD VSS wl[283] BL BLB sram_6t
x_cell284 VDD VSS wl[284] BL BLB sram_6t
x_cell285 VDD VSS wl[285] BL BLB sram_6t
x_cell286 VDD VSS wl[286] BL BLB sram_6t
x_cell287 VDD VSS wl[287] BL BLB sram_6t
x_cell288 VDD VSS wl[288] BL BLB sram_6t
x_cell289 VDD VSS wl[289] BL BLB sram_6t
x_cell290 VDD VSS wl[290] BL BLB sram_6t
x_cell291 VDD VSS wl[291] BL BLB sram_6t
x_cell292 VDD VSS wl[292] BL BLB sram_6t
x_cell293 VDD VSS wl[293] BL BLB sram_6t
x_cell294 VDD VSS wl[294] BL BLB sram_6t
x_cell295 VDD VSS wl[295] BL BLB sram_6t
x_cell296 VDD VSS wl[296] BL BLB sram_6t
x_cell297 VDD VSS wl[297] BL BLB sram_6t
x_cell298 VDD VSS wl[298] BL BLB sram_6t
x_cell299 VDD VSS wl[299] BL BLB sram_6t
x_cell300 VDD VSS wl[300] BL BLB sram_6t
x_cell301 VDD VSS wl[301] BL BLB sram_6t
x_cell302 VDD VSS wl[302] BL BLB sram_6t
x_cell303 VDD VSS wl[303] BL BLB sram_6t
x_cell304 VDD VSS wl[304] BL BLB sram_6t
x_cell305 VDD VSS wl[305] BL BLB sram_6t
x_cell306 VDD VSS wl[306] BL BLB sram_6t
x_cell307 VDD VSS wl[307] BL BLB sram_6t
x_cell308 VDD VSS wl[308] BL BLB sram_6t
x_cell309 VDD VSS wl[309] BL BLB sram_6t
x_cell310 VDD VSS wl[310] BL BLB sram_6t
x_cell311 VDD VSS wl[311] BL BLB sram_6t
x_cell312 VDD VSS wl[312] BL BLB sram_6t
x_cell313 VDD VSS wl[313] BL BLB sram_6t
x_cell314 VDD VSS wl[314] BL BLB sram_6t
x_cell315 VDD VSS wl[315] BL BLB sram_6t
x_cell316 VDD VSS wl[316] BL BLB sram_6t
x_cell317 VDD VSS wl[317] BL BLB sram_6t
x_cell318 VDD VSS wl[318] BL BLB sram_6t
x_cell319 VDD VSS wl[319] BL BLB sram_6t
x_cell320 VDD VSS wl[320] BL BLB sram_6t
x_cell321 VDD VSS wl[321] BL BLB sram_6t
x_cell322 VDD VSS wl[322] BL BLB sram_6t
x_cell323 VDD VSS wl[323] BL BLB sram_6t
x_cell324 VDD VSS wl[324] BL BLB sram_6t
x_cell325 VDD VSS wl[325] BL BLB sram_6t
x_cell326 VDD VSS wl[326] BL BLB sram_6t
x_cell327 VDD VSS wl[327] BL BLB sram_6t
x_cell328 VDD VSS wl[328] BL BLB sram_6t
x_cell329 VDD VSS wl[329] BL BLB sram_6t
x_cell330 VDD VSS wl[330] BL BLB sram_6t
x_cell331 VDD VSS wl[331] BL BLB sram_6t
x_cell332 VDD VSS wl[332] BL BLB sram_6t
x_cell333 VDD VSS wl[333] BL BLB sram_6t
x_cell334 VDD VSS wl[334] BL BLB sram_6t
x_cell335 VDD VSS wl[335] BL BLB sram_6t
x_cell336 VDD VSS wl[336] BL BLB sram_6t
x_cell337 VDD VSS wl[337] BL BLB sram_6t
x_cell338 VDD VSS wl[338] BL BLB sram_6t
x_cell339 VDD VSS wl[339] BL BLB sram_6t
x_cell340 VDD VSS wl[340] BL BLB sram_6t
x_cell341 VDD VSS wl[341] BL BLB sram_6t
x_cell342 VDD VSS wl[342] BL BLB sram_6t
x_cell343 VDD VSS wl[343] BL BLB sram_6t
x_cell344 VDD VSS wl[344] BL BLB sram_6t
x_cell345 VDD VSS wl[345] BL BLB sram_6t
x_cell346 VDD VSS wl[346] BL BLB sram_6t
x_cell347 VDD VSS wl[347] BL BLB sram_6t
x_cell348 VDD VSS wl[348] BL BLB sram_6t
x_cell349 VDD VSS wl[349] BL BLB sram_6t
x_cell350 VDD VSS wl[350] BL BLB sram_6t
x_cell351 VDD VSS wl[351] BL BLB sram_6t
x_cell352 VDD VSS wl[352] BL BLB sram_6t
x_cell353 VDD VSS wl[353] BL BLB sram_6t
x_cell354 VDD VSS wl[354] BL BLB sram_6t
x_cell355 VDD VSS wl[355] BL BLB sram_6t
x_cell356 VDD VSS wl[356] BL BLB sram_6t
x_cell357 VDD VSS wl[357] BL BLB sram_6t
x_cell358 VDD VSS wl[358] BL BLB sram_6t
x_cell359 VDD VSS wl[359] BL BLB sram_6t
x_cell360 VDD VSS wl[360] BL BLB sram_6t
x_cell361 VDD VSS wl[361] BL BLB sram_6t
x_cell362 VDD VSS wl[362] BL BLB sram_6t
x_cell363 VDD VSS wl[363] BL BLB sram_6t
x_cell364 VDD VSS wl[364] BL BLB sram_6t
x_cell365 VDD VSS wl[365] BL BLB sram_6t
x_cell366 VDD VSS wl[366] BL BLB sram_6t
x_cell367 VDD VSS wl[367] BL BLB sram_6t
x_cell368 VDD VSS wl[368] BL BLB sram_6t
x_cell369 VDD VSS wl[369] BL BLB sram_6t
x_cell370 VDD VSS wl[370] BL BLB sram_6t
x_cell371 VDD VSS wl[371] BL BLB sram_6t
x_cell372 VDD VSS wl[372] BL BLB sram_6t
x_cell373 VDD VSS wl[373] BL BLB sram_6t
x_cell374 VDD VSS wl[374] BL BLB sram_6t
x_cell375 VDD VSS wl[375] BL BLB sram_6t
x_cell376 VDD VSS wl[376] BL BLB sram_6t
x_cell377 VDD VSS wl[377] BL BLB sram_6t
x_cell378 VDD VSS wl[378] BL BLB sram_6t
x_cell379 VDD VSS wl[379] BL BLB sram_6t
x_cell380 VDD VSS wl[380] BL BLB sram_6t
x_cell381 VDD VSS wl[381] BL BLB sram_6t
x_cell382 VDD VSS wl[382] BL BLB sram_6t
x_cell383 VDD VSS wl[383] BL BLB sram_6t
x_cell384 VDD VSS wl[384] BL BLB sram_6t
x_cell385 VDD VSS wl[385] BL BLB sram_6t
x_cell386 VDD VSS wl[386] BL BLB sram_6t
x_cell387 VDD VSS wl[387] BL BLB sram_6t
x_cell388 VDD VSS wl[388] BL BLB sram_6t
x_cell389 VDD VSS wl[389] BL BLB sram_6t
x_cell390 VDD VSS wl[390] BL BLB sram_6t
x_cell391 VDD VSS wl[391] BL BLB sram_6t
x_cell392 VDD VSS wl[392] BL BLB sram_6t
x_cell393 VDD VSS wl[393] BL BLB sram_6t
x_cell394 VDD VSS wl[394] BL BLB sram_6t
x_cell395 VDD VSS wl[395] BL BLB sram_6t
x_cell396 VDD VSS wl[396] BL BLB sram_6t
x_cell397 VDD VSS wl[397] BL BLB sram_6t
x_cell398 VDD VSS wl[398] BL BLB sram_6t
x_cell399 VDD VSS wl[399] BL BLB sram_6t
x_cell400 VDD VSS wl[400] BL BLB sram_6t
x_cell401 VDD VSS wl[401] BL BLB sram_6t
x_cell402 VDD VSS wl[402] BL BLB sram_6t
x_cell403 VDD VSS wl[403] BL BLB sram_6t
x_cell404 VDD VSS wl[404] BL BLB sram_6t
x_cell405 VDD VSS wl[405] BL BLB sram_6t
x_cell406 VDD VSS wl[406] BL BLB sram_6t
x_cell407 VDD VSS wl[407] BL BLB sram_6t
x_cell408 VDD VSS wl[408] BL BLB sram_6t
x_cell409 VDD VSS wl[409] BL BLB sram_6t
x_cell410 VDD VSS wl[410] BL BLB sram_6t
x_cell411 VDD VSS wl[411] BL BLB sram_6t
x_cell412 VDD VSS wl[412] BL BLB sram_6t
x_cell413 VDD VSS wl[413] BL BLB sram_6t
x_cell414 VDD VSS wl[414] BL BLB sram_6t
x_cell415 VDD VSS wl[415] BL BLB sram_6t
x_cell416 VDD VSS wl[416] BL BLB sram_6t
x_cell417 VDD VSS wl[417] BL BLB sram_6t
x_cell418 VDD VSS wl[418] BL BLB sram_6t
x_cell419 VDD VSS wl[419] BL BLB sram_6t
x_cell420 VDD VSS wl[420] BL BLB sram_6t
x_cell421 VDD VSS wl[421] BL BLB sram_6t
x_cell422 VDD VSS wl[422] BL BLB sram_6t
x_cell423 VDD VSS wl[423] BL BLB sram_6t
x_cell424 VDD VSS wl[424] BL BLB sram_6t
x_cell425 VDD VSS wl[425] BL BLB sram_6t
x_cell426 VDD VSS wl[426] BL BLB sram_6t
x_cell427 VDD VSS wl[427] BL BLB sram_6t
x_cell428 VDD VSS wl[428] BL BLB sram_6t
x_cell429 VDD VSS wl[429] BL BLB sram_6t
x_cell430 VDD VSS wl[430] BL BLB sram_6t
x_cell431 VDD VSS wl[431] BL BLB sram_6t
x_cell432 VDD VSS wl[432] BL BLB sram_6t
x_cell433 VDD VSS wl[433] BL BLB sram_6t
x_cell434 VDD VSS wl[434] BL BLB sram_6t
x_cell435 VDD VSS wl[435] BL BLB sram_6t
x_cell436 VDD VSS wl[436] BL BLB sram_6t
x_cell437 VDD VSS wl[437] BL BLB sram_6t
x_cell438 VDD VSS wl[438] BL BLB sram_6t
x_cell439 VDD VSS wl[439] BL BLB sram_6t
x_cell440 VDD VSS wl[440] BL BLB sram_6t
x_cell441 VDD VSS wl[441] BL BLB sram_6t
x_cell442 VDD VSS wl[442] BL BLB sram_6t
x_cell443 VDD VSS wl[443] BL BLB sram_6t
x_cell444 VDD VSS wl[444] BL BLB sram_6t
x_cell445 VDD VSS wl[445] BL BLB sram_6t
x_cell446 VDD VSS wl[446] BL BLB sram_6t
x_cell447 VDD VSS wl[447] BL BLB sram_6t
x_cell448 VDD VSS wl[448] BL BLB sram_6t
x_cell449 VDD VSS wl[449] BL BLB sram_6t
x_cell450 VDD VSS wl[450] BL BLB sram_6t
x_cell451 VDD VSS wl[451] BL BLB sram_6t
x_cell452 VDD VSS wl[452] BL BLB sram_6t
x_cell453 VDD VSS wl[453] BL BLB sram_6t
x_cell454 VDD VSS wl[454] BL BLB sram_6t
x_cell455 VDD VSS wl[455] BL BLB sram_6t
x_cell456 VDD VSS wl[456] BL BLB sram_6t
x_cell457 VDD VSS wl[457] BL BLB sram_6t
x_cell458 VDD VSS wl[458] BL BLB sram_6t
x_cell459 VDD VSS wl[459] BL BLB sram_6t
x_cell460 VDD VSS wl[460] BL BLB sram_6t
x_cell461 VDD VSS wl[461] BL BLB sram_6t
x_cell462 VDD VSS wl[462] BL BLB sram_6t
x_cell463 VDD VSS wl[463] BL BLB sram_6t
x_cell464 VDD VSS wl[464] BL BLB sram_6t
x_cell465 VDD VSS wl[465] BL BLB sram_6t
x_cell466 VDD VSS wl[466] BL BLB sram_6t
x_cell467 VDD VSS wl[467] BL BLB sram_6t
x_cell468 VDD VSS wl[468] BL BLB sram_6t
x_cell469 VDD VSS wl[469] BL BLB sram_6t
x_cell470 VDD VSS wl[470] BL BLB sram_6t
x_cell471 VDD VSS wl[471] BL BLB sram_6t
x_cell472 VDD VSS wl[472] BL BLB sram_6t
x_cell473 VDD VSS wl[473] BL BLB sram_6t
x_cell474 VDD VSS wl[474] BL BLB sram_6t
x_cell475 VDD VSS wl[475] BL BLB sram_6t
x_cell476 VDD VSS wl[476] BL BLB sram_6t
x_cell477 VDD VSS wl[477] BL BLB sram_6t
x_cell478 VDD VSS wl[478] BL BLB sram_6t
x_cell479 VDD VSS wl[479] BL BLB sram_6t
x_cell480 VDD VSS wl[480] BL BLB sram_6t
x_cell481 VDD VSS wl[481] BL BLB sram_6t
x_cell482 VDD VSS wl[482] BL BLB sram_6t
x_cell483 VDD VSS wl[483] BL BLB sram_6t
x_cell484 VDD VSS wl[484] BL BLB sram_6t
x_cell485 VDD VSS wl[485] BL BLB sram_6t
x_cell486 VDD VSS wl[486] BL BLB sram_6t
x_cell487 VDD VSS wl[487] BL BLB sram_6t
x_cell488 VDD VSS wl[488] BL BLB sram_6t
x_cell489 VDD VSS wl[489] BL BLB sram_6t
x_cell490 VDD VSS wl[490] BL BLB sram_6t
x_cell491 VDD VSS wl[491] BL BLB sram_6t
x_cell492 VDD VSS wl[492] BL BLB sram_6t
x_cell493 VDD VSS wl[493] BL BLB sram_6t
x_cell494 VDD VSS wl[494] BL BLB sram_6t
x_cell495 VDD VSS wl[495] BL BLB sram_6t
x_cell496 VDD VSS wl[496] BL BLB sram_6t
x_cell497 VDD VSS wl[497] BL BLB sram_6t
x_cell498 VDD VSS wl[498] BL BLB sram_6t
x_cell499 VDD VSS wl[499] BL BLB sram_6t
x_cell500 VDD VSS wl[500] BL BLB sram_6t
x_cell501 VDD VSS wl[501] BL BLB sram_6t
x_cell502 VDD VSS wl[502] BL BLB sram_6t
x_cell503 VDD VSS wl[503] BL BLB sram_6t
x_cell504 VDD VSS wl[504] BL BLB sram_6t
x_cell505 VDD VSS wl[505] BL BLB sram_6t
x_cell506 VDD VSS wl[506] BL BLB sram_6t
x_cell507 VDD VSS wl[507] BL BLB sram_6t
x_cell508 VDD VSS wl[508] BL BLB sram_6t
x_cell509 VDD VSS wl[509] BL BLB sram_6t
x_cell510 VDD VSS wl[510] BL BLB sram_6t
x_cell511 VDD VSS wl[511] BL BLB sram_6t
.ends
.subckt buffer_arr512 VDD VSS clk
+ in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7]
+ in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15]
+ in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23]
+ in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31]
+ in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39]
+ in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47]
+ in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55]
+ in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63]
+ in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71]
+ in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79]
+ in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87]
+ in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95]
+ in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103]
+ in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111]
+ in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119]
+ in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127]
+ in[128] in[129] in[130] in[131] in[132] in[133] in[134] in[135]
+ in[136] in[137] in[138] in[139] in[140] in[141] in[142] in[143]
+ in[144] in[145] in[146] in[147] in[148] in[149] in[150] in[151]
+ in[152] in[153] in[154] in[155] in[156] in[157] in[158] in[159]
+ in[160] in[161] in[162] in[163] in[164] in[165] in[166] in[167]
+ in[168] in[169] in[170] in[171] in[172] in[173] in[174] in[175]
+ in[176] in[177] in[178] in[179] in[180] in[181] in[182] in[183]
+ in[184] in[185] in[186] in[187] in[188] in[189] in[190] in[191]
+ in[192] in[193] in[194] in[195] in[196] in[197] in[198] in[199]
+ in[200] in[201] in[202] in[203] in[204] in[205] in[206] in[207]
+ in[208] in[209] in[210] in[211] in[212] in[213] in[214] in[215]
+ in[216] in[217] in[218] in[219] in[220] in[221] in[222] in[223]
+ in[224] in[225] in[226] in[227] in[228] in[229] in[230] in[231]
+ in[232] in[233] in[234] in[235] in[236] in[237] in[238] in[239]
+ in[240] in[241] in[242] in[243] in[244] in[245] in[246] in[247]
+ in[248] in[249] in[250] in[251] in[252] in[253] in[254] in[255]
+ in[256] in[257] in[258] in[259] in[260] in[261] in[262] in[263]
+ in[264] in[265] in[266] in[267] in[268] in[269] in[270] in[271]
+ in[272] in[273] in[274] in[275] in[276] in[277] in[278] in[279]
+ in[280] in[281] in[282] in[283] in[284] in[285] in[286] in[287]
+ in[288] in[289] in[290] in[291] in[292] in[293] in[294] in[295]
+ in[296] in[297] in[298] in[299] in[300] in[301] in[302] in[303]
+ in[304] in[305] in[306] in[307] in[308] in[309] in[310] in[311]
+ in[312] in[313] in[314] in[315] in[316] in[317] in[318] in[319]
+ in[320] in[321] in[322] in[323] in[324] in[325] in[326] in[327]
+ in[328] in[329] in[330] in[331] in[332] in[333] in[334] in[335]
+ in[336] in[337] in[338] in[339] in[340] in[341] in[342] in[343]
+ in[344] in[345] in[346] in[347] in[348] in[349] in[350] in[351]
+ in[352] in[353] in[354] in[355] in[356] in[357] in[358] in[359]
+ in[360] in[361] in[362] in[363] in[364] in[365] in[366] in[367]
+ in[368] in[369] in[370] in[371] in[372] in[373] in[374] in[375]
+ in[376] in[377] in[378] in[379] in[380] in[381] in[382] in[383]
+ in[384] in[385] in[386] in[387] in[388] in[389] in[390] in[391]
+ in[392] in[393] in[394] in[395] in[396] in[397] in[398] in[399]
+ in[400] in[401] in[402] in[403] in[404] in[405] in[406] in[407]
+ in[408] in[409] in[410] in[411] in[412] in[413] in[414] in[415]
+ in[416] in[417] in[418] in[419] in[420] in[421] in[422] in[423]
+ in[424] in[425] in[426] in[427] in[428] in[429] in[430] in[431]
+ in[432] in[433] in[434] in[435] in[436] in[437] in[438] in[439]
+ in[440] in[441] in[442] in[443] in[444] in[445] in[446] in[447]
+ in[448] in[449] in[450] in[451] in[452] in[453] in[454] in[455]
+ in[456] in[457] in[458] in[459] in[460] in[461] in[462] in[463]
+ in[464] in[465] in[466] in[467] in[468] in[469] in[470] in[471]
+ in[472] in[473] in[474] in[475] in[476] in[477] in[478] in[479]
+ in[480] in[481] in[482] in[483] in[484] in[485] in[486] in[487]
+ in[488] in[489] in[490] in[491] in[492] in[493] in[494] in[495]
+ in[496] in[497] in[498] in[499] in[500] in[501] in[502] in[503]
+ in[504] in[505] in[506] in[507] in[508] in[509] in[510] in[511]
+ out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7]
+ out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15]
+ out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23]
+ out[24] out[25] out[26] out[27] out[28] out[29] out[30] out[31]
+ out[32] out[33] out[34] out[35] out[36] out[37] out[38] out[39]
+ out[40] out[41] out[42] out[43] out[44] out[45] out[46] out[47]
+ out[48] out[49] out[50] out[51] out[52] out[53] out[54] out[55]
+ out[56] out[57] out[58] out[59] out[60] out[61] out[62] out[63]
+ out[64] out[65] out[66] out[67] out[68] out[69] out[70] out[71]
+ out[72] out[73] out[74] out[75] out[76] out[77] out[78] out[79]
+ out[80] out[81] out[82] out[83] out[84] out[85] out[86] out[87]
+ out[88] out[89] out[90] out[91] out[92] out[93] out[94] out[95]
+ out[96] out[97] out[98] out[99] out[100] out[101] out[102] out[103]
+ out[104] out[105] out[106] out[107] out[108] out[109] out[110] out[111]
+ out[112] out[113] out[114] out[115] out[116] out[117] out[118] out[119]
+ out[120] out[121] out[122] out[123] out[124] out[125] out[126] out[127]
+ out[128] out[129] out[130] out[131] out[132] out[133] out[134] out[135]
+ out[136] out[137] out[138] out[139] out[140] out[141] out[142] out[143]
+ out[144] out[145] out[146] out[147] out[148] out[149] out[150] out[151]
+ out[152] out[153] out[154] out[155] out[156] out[157] out[158] out[159]
+ out[160] out[161] out[162] out[163] out[164] out[165] out[166] out[167]
+ out[168] out[169] out[170] out[171] out[172] out[173] out[174] out[175]
+ out[176] out[177] out[178] out[179] out[180] out[181] out[182] out[183]
+ out[184] out[185] out[186] out[187] out[188] out[189] out[190] out[191]
+ out[192] out[193] out[194] out[195] out[196] out[197] out[198] out[199]
+ out[200] out[201] out[202] out[203] out[204] out[205] out[206] out[207]
+ out[208] out[209] out[210] out[211] out[212] out[213] out[214] out[215]
+ out[216] out[217] out[218] out[219] out[220] out[221] out[222] out[223]
+ out[224] out[225] out[226] out[227] out[228] out[229] out[230] out[231]
+ out[232] out[233] out[234] out[235] out[236] out[237] out[238] out[239]
+ out[240] out[241] out[242] out[243] out[244] out[245] out[246] out[247]
+ out[248] out[249] out[250] out[251] out[252] out[253] out[254] out[255]
+ out[256] out[257] out[258] out[259] out[260] out[261] out[262] out[263]
+ out[264] out[265] out[266] out[267] out[268] out[269] out[270] out[271]
+ out[272] out[273] out[274] out[275] out[276] out[277] out[278] out[279]
+ out[280] out[281] out[282] out[283] out[284] out[285] out[286] out[287]
+ out[288] out[289] out[290] out[291] out[292] out[293] out[294] out[295]
+ out[296] out[297] out[298] out[299] out[300] out[301] out[302] out[303]
+ out[304] out[305] out[306] out[307] out[308] out[309] out[310] out[311]
+ out[312] out[313] out[314] out[315] out[316] out[317] out[318] out[319]
+ out[320] out[321] out[322] out[323] out[324] out[325] out[326] out[327]
+ out[328] out[329] out[330] out[331] out[332] out[333] out[334] out[335]
+ out[336] out[337] out[338] out[339] out[340] out[341] out[342] out[343]
+ out[344] out[345] out[346] out[347] out[348] out[349] out[350] out[351]
+ out[352] out[353] out[354] out[355] out[356] out[357] out[358] out[359]
+ out[360] out[361] out[362] out[363] out[364] out[365] out[366] out[367]
+ out[368] out[369] out[370] out[371] out[372] out[373] out[374] out[375]
+ out[376] out[377] out[378] out[379] out[380] out[381] out[382] out[383]
+ out[384] out[385] out[386] out[387] out[388] out[389] out[390] out[391]
+ out[392] out[393] out[394] out[395] out[396] out[397] out[398] out[399]
+ out[400] out[401] out[402] out[403] out[404] out[405] out[406] out[407]
+ out[408] out[409] out[410] out[411] out[412] out[413] out[414] out[415]
+ out[416] out[417] out[418] out[419] out[420] out[421] out[422] out[423]
+ out[424] out[425] out[426] out[427] out[428] out[429] out[430] out[431]
+ out[432] out[433] out[434] out[435] out[436] out[437] out[438] out[439]
+ out[440] out[441] out[442] out[443] out[444] out[445] out[446] out[447]
+ out[448] out[449] out[450] out[451] out[452] out[453] out[454] out[455]
+ out[456] out[457] out[458] out[459] out[460] out[461] out[462] out[463]
+ out[464] out[465] out[466] out[467] out[468] out[469] out[470] out[471]
+ out[472] out[473] out[474] out[475] out[476] out[477] out[478] out[479]
+ out[480] out[481] out[482] out[483] out[484] out[485] out[486] out[487]
+ out[488] out[489] out[490] out[491] out[492] out[493] out[494] out[495]
+ out[496] out[497] out[498] out[499] out[500] out[501] out[502] out[503]
+ out[504] out[505] out[506] out[507] out[508] out[509] out[510] out[511]
x_buf0 VDD VSS in[0] out[0] buffer
x_and0 VSS VDD in[0] clk out[0] AND2x2_ASAP7_75t_SRAM
x_buf1 VDD VSS in[1] out[1] buffer
x_and1 VSS VDD in[1] clk out[1] AND2x2_ASAP7_75t_SRAM
x_buf2 VDD VSS in[2] out[2] buffer
x_and2 VSS VDD in[2] clk out[2] AND2x2_ASAP7_75t_SRAM
x_buf3 VDD VSS in[3] out[3] buffer
x_and3 VSS VDD in[3] clk out[3] AND2x2_ASAP7_75t_SRAM
x_buf4 VDD VSS in[4] out[4] buffer
x_and4 VSS VDD in[4] clk out[4] AND2x2_ASAP7_75t_SRAM
x_buf5 VDD VSS in[5] out[5] buffer
x_and5 VSS VDD in[5] clk out[5] AND2x2_ASAP7_75t_SRAM
x_buf6 VDD VSS in[6] out[6] buffer
x_and6 VSS VDD in[6] clk out[6] AND2x2_ASAP7_75t_SRAM
x_buf7 VDD VSS in[7] out[7] buffer
x_and7 VSS VDD in[7] clk out[7] AND2x2_ASAP7_75t_SRAM
x_buf8 VDD VSS in[8] out[8] buffer
x_and8 VSS VDD in[8] clk out[8] AND2x2_ASAP7_75t_SRAM
x_buf9 VDD VSS in[9] out[9] buffer
x_and9 VSS VDD in[9] clk out[9] AND2x2_ASAP7_75t_SRAM
x_buf10 VDD VSS in[10] out[10] buffer
x_and10 VSS VDD in[10] clk out[10] AND2x2_ASAP7_75t_SRAM
x_buf11 VDD VSS in[11] out[11] buffer
x_and11 VSS VDD in[11] clk out[11] AND2x2_ASAP7_75t_SRAM
x_buf12 VDD VSS in[12] out[12] buffer
x_and12 VSS VDD in[12] clk out[12] AND2x2_ASAP7_75t_SRAM
x_buf13 VDD VSS in[13] out[13] buffer
x_and13 VSS VDD in[13] clk out[13] AND2x2_ASAP7_75t_SRAM
x_buf14 VDD VSS in[14] out[14] buffer
x_and14 VSS VDD in[14] clk out[14] AND2x2_ASAP7_75t_SRAM
x_buf15 VDD VSS in[15] out[15] buffer
x_and15 VSS VDD in[15] clk out[15] AND2x2_ASAP7_75t_SRAM
x_buf16 VDD VSS in[16] out[16] buffer
x_and16 VSS VDD in[16] clk out[16] AND2x2_ASAP7_75t_SRAM
x_buf17 VDD VSS in[17] out[17] buffer
x_and17 VSS VDD in[17] clk out[17] AND2x2_ASAP7_75t_SRAM
x_buf18 VDD VSS in[18] out[18] buffer
x_and18 VSS VDD in[18] clk out[18] AND2x2_ASAP7_75t_SRAM
x_buf19 VDD VSS in[19] out[19] buffer
x_and19 VSS VDD in[19] clk out[19] AND2x2_ASAP7_75t_SRAM
x_buf20 VDD VSS in[20] out[20] buffer
x_and20 VSS VDD in[20] clk out[20] AND2x2_ASAP7_75t_SRAM
x_buf21 VDD VSS in[21] out[21] buffer
x_and21 VSS VDD in[21] clk out[21] AND2x2_ASAP7_75t_SRAM
x_buf22 VDD VSS in[22] out[22] buffer
x_and22 VSS VDD in[22] clk out[22] AND2x2_ASAP7_75t_SRAM
x_buf23 VDD VSS in[23] out[23] buffer
x_and23 VSS VDD in[23] clk out[23] AND2x2_ASAP7_75t_SRAM
x_buf24 VDD VSS in[24] out[24] buffer
x_and24 VSS VDD in[24] clk out[24] AND2x2_ASAP7_75t_SRAM
x_buf25 VDD VSS in[25] out[25] buffer
x_and25 VSS VDD in[25] clk out[25] AND2x2_ASAP7_75t_SRAM
x_buf26 VDD VSS in[26] out[26] buffer
x_and26 VSS VDD in[26] clk out[26] AND2x2_ASAP7_75t_SRAM
x_buf27 VDD VSS in[27] out[27] buffer
x_and27 VSS VDD in[27] clk out[27] AND2x2_ASAP7_75t_SRAM
x_buf28 VDD VSS in[28] out[28] buffer
x_and28 VSS VDD in[28] clk out[28] AND2x2_ASAP7_75t_SRAM
x_buf29 VDD VSS in[29] out[29] buffer
x_and29 VSS VDD in[29] clk out[29] AND2x2_ASAP7_75t_SRAM
x_buf30 VDD VSS in[30] out[30] buffer
x_and30 VSS VDD in[30] clk out[30] AND2x2_ASAP7_75t_SRAM
x_buf31 VDD VSS in[31] out[31] buffer
x_and31 VSS VDD in[31] clk out[31] AND2x2_ASAP7_75t_SRAM
x_buf32 VDD VSS in[32] out[32] buffer
x_and32 VSS VDD in[32] clk out[32] AND2x2_ASAP7_75t_SRAM
x_buf33 VDD VSS in[33] out[33] buffer
x_and33 VSS VDD in[33] clk out[33] AND2x2_ASAP7_75t_SRAM
x_buf34 VDD VSS in[34] out[34] buffer
x_and34 VSS VDD in[34] clk out[34] AND2x2_ASAP7_75t_SRAM
x_buf35 VDD VSS in[35] out[35] buffer
x_and35 VSS VDD in[35] clk out[35] AND2x2_ASAP7_75t_SRAM
x_buf36 VDD VSS in[36] out[36] buffer
x_and36 VSS VDD in[36] clk out[36] AND2x2_ASAP7_75t_SRAM
x_buf37 VDD VSS in[37] out[37] buffer
x_and37 VSS VDD in[37] clk out[37] AND2x2_ASAP7_75t_SRAM
x_buf38 VDD VSS in[38] out[38] buffer
x_and38 VSS VDD in[38] clk out[38] AND2x2_ASAP7_75t_SRAM
x_buf39 VDD VSS in[39] out[39] buffer
x_and39 VSS VDD in[39] clk out[39] AND2x2_ASAP7_75t_SRAM
x_buf40 VDD VSS in[40] out[40] buffer
x_and40 VSS VDD in[40] clk out[40] AND2x2_ASAP7_75t_SRAM
x_buf41 VDD VSS in[41] out[41] buffer
x_and41 VSS VDD in[41] clk out[41] AND2x2_ASAP7_75t_SRAM
x_buf42 VDD VSS in[42] out[42] buffer
x_and42 VSS VDD in[42] clk out[42] AND2x2_ASAP7_75t_SRAM
x_buf43 VDD VSS in[43] out[43] buffer
x_and43 VSS VDD in[43] clk out[43] AND2x2_ASAP7_75t_SRAM
x_buf44 VDD VSS in[44] out[44] buffer
x_and44 VSS VDD in[44] clk out[44] AND2x2_ASAP7_75t_SRAM
x_buf45 VDD VSS in[45] out[45] buffer
x_and45 VSS VDD in[45] clk out[45] AND2x2_ASAP7_75t_SRAM
x_buf46 VDD VSS in[46] out[46] buffer
x_and46 VSS VDD in[46] clk out[46] AND2x2_ASAP7_75t_SRAM
x_buf47 VDD VSS in[47] out[47] buffer
x_and47 VSS VDD in[47] clk out[47] AND2x2_ASAP7_75t_SRAM
x_buf48 VDD VSS in[48] out[48] buffer
x_and48 VSS VDD in[48] clk out[48] AND2x2_ASAP7_75t_SRAM
x_buf49 VDD VSS in[49] out[49] buffer
x_and49 VSS VDD in[49] clk out[49] AND2x2_ASAP7_75t_SRAM
x_buf50 VDD VSS in[50] out[50] buffer
x_and50 VSS VDD in[50] clk out[50] AND2x2_ASAP7_75t_SRAM
x_buf51 VDD VSS in[51] out[51] buffer
x_and51 VSS VDD in[51] clk out[51] AND2x2_ASAP7_75t_SRAM
x_buf52 VDD VSS in[52] out[52] buffer
x_and52 VSS VDD in[52] clk out[52] AND2x2_ASAP7_75t_SRAM
x_buf53 VDD VSS in[53] out[53] buffer
x_and53 VSS VDD in[53] clk out[53] AND2x2_ASAP7_75t_SRAM
x_buf54 VDD VSS in[54] out[54] buffer
x_and54 VSS VDD in[54] clk out[54] AND2x2_ASAP7_75t_SRAM
x_buf55 VDD VSS in[55] out[55] buffer
x_and55 VSS VDD in[55] clk out[55] AND2x2_ASAP7_75t_SRAM
x_buf56 VDD VSS in[56] out[56] buffer
x_and56 VSS VDD in[56] clk out[56] AND2x2_ASAP7_75t_SRAM
x_buf57 VDD VSS in[57] out[57] buffer
x_and57 VSS VDD in[57] clk out[57] AND2x2_ASAP7_75t_SRAM
x_buf58 VDD VSS in[58] out[58] buffer
x_and58 VSS VDD in[58] clk out[58] AND2x2_ASAP7_75t_SRAM
x_buf59 VDD VSS in[59] out[59] buffer
x_and59 VSS VDD in[59] clk out[59] AND2x2_ASAP7_75t_SRAM
x_buf60 VDD VSS in[60] out[60] buffer
x_and60 VSS VDD in[60] clk out[60] AND2x2_ASAP7_75t_SRAM
x_buf61 VDD VSS in[61] out[61] buffer
x_and61 VSS VDD in[61] clk out[61] AND2x2_ASAP7_75t_SRAM
x_buf62 VDD VSS in[62] out[62] buffer
x_and62 VSS VDD in[62] clk out[62] AND2x2_ASAP7_75t_SRAM
x_buf63 VDD VSS in[63] out[63] buffer
x_and63 VSS VDD in[63] clk out[63] AND2x2_ASAP7_75t_SRAM
x_buf64 VDD VSS in[64] out[64] buffer
x_and64 VSS VDD in[64] clk out[64] AND2x2_ASAP7_75t_SRAM
x_buf65 VDD VSS in[65] out[65] buffer
x_and65 VSS VDD in[65] clk out[65] AND2x2_ASAP7_75t_SRAM
x_buf66 VDD VSS in[66] out[66] buffer
x_and66 VSS VDD in[66] clk out[66] AND2x2_ASAP7_75t_SRAM
x_buf67 VDD VSS in[67] out[67] buffer
x_and67 VSS VDD in[67] clk out[67] AND2x2_ASAP7_75t_SRAM
x_buf68 VDD VSS in[68] out[68] buffer
x_and68 VSS VDD in[68] clk out[68] AND2x2_ASAP7_75t_SRAM
x_buf69 VDD VSS in[69] out[69] buffer
x_and69 VSS VDD in[69] clk out[69] AND2x2_ASAP7_75t_SRAM
x_buf70 VDD VSS in[70] out[70] buffer
x_and70 VSS VDD in[70] clk out[70] AND2x2_ASAP7_75t_SRAM
x_buf71 VDD VSS in[71] out[71] buffer
x_and71 VSS VDD in[71] clk out[71] AND2x2_ASAP7_75t_SRAM
x_buf72 VDD VSS in[72] out[72] buffer
x_and72 VSS VDD in[72] clk out[72] AND2x2_ASAP7_75t_SRAM
x_buf73 VDD VSS in[73] out[73] buffer
x_and73 VSS VDD in[73] clk out[73] AND2x2_ASAP7_75t_SRAM
x_buf74 VDD VSS in[74] out[74] buffer
x_and74 VSS VDD in[74] clk out[74] AND2x2_ASAP7_75t_SRAM
x_buf75 VDD VSS in[75] out[75] buffer
x_and75 VSS VDD in[75] clk out[75] AND2x2_ASAP7_75t_SRAM
x_buf76 VDD VSS in[76] out[76] buffer
x_and76 VSS VDD in[76] clk out[76] AND2x2_ASAP7_75t_SRAM
x_buf77 VDD VSS in[77] out[77] buffer
x_and77 VSS VDD in[77] clk out[77] AND2x2_ASAP7_75t_SRAM
x_buf78 VDD VSS in[78] out[78] buffer
x_and78 VSS VDD in[78] clk out[78] AND2x2_ASAP7_75t_SRAM
x_buf79 VDD VSS in[79] out[79] buffer
x_and79 VSS VDD in[79] clk out[79] AND2x2_ASAP7_75t_SRAM
x_buf80 VDD VSS in[80] out[80] buffer
x_and80 VSS VDD in[80] clk out[80] AND2x2_ASAP7_75t_SRAM
x_buf81 VDD VSS in[81] out[81] buffer
x_and81 VSS VDD in[81] clk out[81] AND2x2_ASAP7_75t_SRAM
x_buf82 VDD VSS in[82] out[82] buffer
x_and82 VSS VDD in[82] clk out[82] AND2x2_ASAP7_75t_SRAM
x_buf83 VDD VSS in[83] out[83] buffer
x_and83 VSS VDD in[83] clk out[83] AND2x2_ASAP7_75t_SRAM
x_buf84 VDD VSS in[84] out[84] buffer
x_and84 VSS VDD in[84] clk out[84] AND2x2_ASAP7_75t_SRAM
x_buf85 VDD VSS in[85] out[85] buffer
x_and85 VSS VDD in[85] clk out[85] AND2x2_ASAP7_75t_SRAM
x_buf86 VDD VSS in[86] out[86] buffer
x_and86 VSS VDD in[86] clk out[86] AND2x2_ASAP7_75t_SRAM
x_buf87 VDD VSS in[87] out[87] buffer
x_and87 VSS VDD in[87] clk out[87] AND2x2_ASAP7_75t_SRAM
x_buf88 VDD VSS in[88] out[88] buffer
x_and88 VSS VDD in[88] clk out[88] AND2x2_ASAP7_75t_SRAM
x_buf89 VDD VSS in[89] out[89] buffer
x_and89 VSS VDD in[89] clk out[89] AND2x2_ASAP7_75t_SRAM
x_buf90 VDD VSS in[90] out[90] buffer
x_and90 VSS VDD in[90] clk out[90] AND2x2_ASAP7_75t_SRAM
x_buf91 VDD VSS in[91] out[91] buffer
x_and91 VSS VDD in[91] clk out[91] AND2x2_ASAP7_75t_SRAM
x_buf92 VDD VSS in[92] out[92] buffer
x_and92 VSS VDD in[92] clk out[92] AND2x2_ASAP7_75t_SRAM
x_buf93 VDD VSS in[93] out[93] buffer
x_and93 VSS VDD in[93] clk out[93] AND2x2_ASAP7_75t_SRAM
x_buf94 VDD VSS in[94] out[94] buffer
x_and94 VSS VDD in[94] clk out[94] AND2x2_ASAP7_75t_SRAM
x_buf95 VDD VSS in[95] out[95] buffer
x_and95 VSS VDD in[95] clk out[95] AND2x2_ASAP7_75t_SRAM
x_buf96 VDD VSS in[96] out[96] buffer
x_and96 VSS VDD in[96] clk out[96] AND2x2_ASAP7_75t_SRAM
x_buf97 VDD VSS in[97] out[97] buffer
x_and97 VSS VDD in[97] clk out[97] AND2x2_ASAP7_75t_SRAM
x_buf98 VDD VSS in[98] out[98] buffer
x_and98 VSS VDD in[98] clk out[98] AND2x2_ASAP7_75t_SRAM
x_buf99 VDD VSS in[99] out[99] buffer
x_and99 VSS VDD in[99] clk out[99] AND2x2_ASAP7_75t_SRAM
x_buf100 VDD VSS in[100] out[100] buffer
x_and100 VSS VDD in[100] clk out[100] AND2x2_ASAP7_75t_SRAM
x_buf101 VDD VSS in[101] out[101] buffer
x_and101 VSS VDD in[101] clk out[101] AND2x2_ASAP7_75t_SRAM
x_buf102 VDD VSS in[102] out[102] buffer
x_and102 VSS VDD in[102] clk out[102] AND2x2_ASAP7_75t_SRAM
x_buf103 VDD VSS in[103] out[103] buffer
x_and103 VSS VDD in[103] clk out[103] AND2x2_ASAP7_75t_SRAM
x_buf104 VDD VSS in[104] out[104] buffer
x_and104 VSS VDD in[104] clk out[104] AND2x2_ASAP7_75t_SRAM
x_buf105 VDD VSS in[105] out[105] buffer
x_and105 VSS VDD in[105] clk out[105] AND2x2_ASAP7_75t_SRAM
x_buf106 VDD VSS in[106] out[106] buffer
x_and106 VSS VDD in[106] clk out[106] AND2x2_ASAP7_75t_SRAM
x_buf107 VDD VSS in[107] out[107] buffer
x_and107 VSS VDD in[107] clk out[107] AND2x2_ASAP7_75t_SRAM
x_buf108 VDD VSS in[108] out[108] buffer
x_and108 VSS VDD in[108] clk out[108] AND2x2_ASAP7_75t_SRAM
x_buf109 VDD VSS in[109] out[109] buffer
x_and109 VSS VDD in[109] clk out[109] AND2x2_ASAP7_75t_SRAM
x_buf110 VDD VSS in[110] out[110] buffer
x_and110 VSS VDD in[110] clk out[110] AND2x2_ASAP7_75t_SRAM
x_buf111 VDD VSS in[111] out[111] buffer
x_and111 VSS VDD in[111] clk out[111] AND2x2_ASAP7_75t_SRAM
x_buf112 VDD VSS in[112] out[112] buffer
x_and112 VSS VDD in[112] clk out[112] AND2x2_ASAP7_75t_SRAM
x_buf113 VDD VSS in[113] out[113] buffer
x_and113 VSS VDD in[113] clk out[113] AND2x2_ASAP7_75t_SRAM
x_buf114 VDD VSS in[114] out[114] buffer
x_and114 VSS VDD in[114] clk out[114] AND2x2_ASAP7_75t_SRAM
x_buf115 VDD VSS in[115] out[115] buffer
x_and115 VSS VDD in[115] clk out[115] AND2x2_ASAP7_75t_SRAM
x_buf116 VDD VSS in[116] out[116] buffer
x_and116 VSS VDD in[116] clk out[116] AND2x2_ASAP7_75t_SRAM
x_buf117 VDD VSS in[117] out[117] buffer
x_and117 VSS VDD in[117] clk out[117] AND2x2_ASAP7_75t_SRAM
x_buf118 VDD VSS in[118] out[118] buffer
x_and118 VSS VDD in[118] clk out[118] AND2x2_ASAP7_75t_SRAM
x_buf119 VDD VSS in[119] out[119] buffer
x_and119 VSS VDD in[119] clk out[119] AND2x2_ASAP7_75t_SRAM
x_buf120 VDD VSS in[120] out[120] buffer
x_and120 VSS VDD in[120] clk out[120] AND2x2_ASAP7_75t_SRAM
x_buf121 VDD VSS in[121] out[121] buffer
x_and121 VSS VDD in[121] clk out[121] AND2x2_ASAP7_75t_SRAM
x_buf122 VDD VSS in[122] out[122] buffer
x_and122 VSS VDD in[122] clk out[122] AND2x2_ASAP7_75t_SRAM
x_buf123 VDD VSS in[123] out[123] buffer
x_and123 VSS VDD in[123] clk out[123] AND2x2_ASAP7_75t_SRAM
x_buf124 VDD VSS in[124] out[124] buffer
x_and124 VSS VDD in[124] clk out[124] AND2x2_ASAP7_75t_SRAM
x_buf125 VDD VSS in[125] out[125] buffer
x_and125 VSS VDD in[125] clk out[125] AND2x2_ASAP7_75t_SRAM
x_buf126 VDD VSS in[126] out[126] buffer
x_and126 VSS VDD in[126] clk out[126] AND2x2_ASAP7_75t_SRAM
x_buf127 VDD VSS in[127] out[127] buffer
x_and127 VSS VDD in[127] clk out[127] AND2x2_ASAP7_75t_SRAM
x_buf128 VDD VSS in[128] out[128] buffer
x_and128 VSS VDD in[128] clk out[128] AND2x2_ASAP7_75t_SRAM
x_buf129 VDD VSS in[129] out[129] buffer
x_and129 VSS VDD in[129] clk out[129] AND2x2_ASAP7_75t_SRAM
x_buf130 VDD VSS in[130] out[130] buffer
x_and130 VSS VDD in[130] clk out[130] AND2x2_ASAP7_75t_SRAM
x_buf131 VDD VSS in[131] out[131] buffer
x_and131 VSS VDD in[131] clk out[131] AND2x2_ASAP7_75t_SRAM
x_buf132 VDD VSS in[132] out[132] buffer
x_and132 VSS VDD in[132] clk out[132] AND2x2_ASAP7_75t_SRAM
x_buf133 VDD VSS in[133] out[133] buffer
x_and133 VSS VDD in[133] clk out[133] AND2x2_ASAP7_75t_SRAM
x_buf134 VDD VSS in[134] out[134] buffer
x_and134 VSS VDD in[134] clk out[134] AND2x2_ASAP7_75t_SRAM
x_buf135 VDD VSS in[135] out[135] buffer
x_and135 VSS VDD in[135] clk out[135] AND2x2_ASAP7_75t_SRAM
x_buf136 VDD VSS in[136] out[136] buffer
x_and136 VSS VDD in[136] clk out[136] AND2x2_ASAP7_75t_SRAM
x_buf137 VDD VSS in[137] out[137] buffer
x_and137 VSS VDD in[137] clk out[137] AND2x2_ASAP7_75t_SRAM
x_buf138 VDD VSS in[138] out[138] buffer
x_and138 VSS VDD in[138] clk out[138] AND2x2_ASAP7_75t_SRAM
x_buf139 VDD VSS in[139] out[139] buffer
x_and139 VSS VDD in[139] clk out[139] AND2x2_ASAP7_75t_SRAM
x_buf140 VDD VSS in[140] out[140] buffer
x_and140 VSS VDD in[140] clk out[140] AND2x2_ASAP7_75t_SRAM
x_buf141 VDD VSS in[141] out[141] buffer
x_and141 VSS VDD in[141] clk out[141] AND2x2_ASAP7_75t_SRAM
x_buf142 VDD VSS in[142] out[142] buffer
x_and142 VSS VDD in[142] clk out[142] AND2x2_ASAP7_75t_SRAM
x_buf143 VDD VSS in[143] out[143] buffer
x_and143 VSS VDD in[143] clk out[143] AND2x2_ASAP7_75t_SRAM
x_buf144 VDD VSS in[144] out[144] buffer
x_and144 VSS VDD in[144] clk out[144] AND2x2_ASAP7_75t_SRAM
x_buf145 VDD VSS in[145] out[145] buffer
x_and145 VSS VDD in[145] clk out[145] AND2x2_ASAP7_75t_SRAM
x_buf146 VDD VSS in[146] out[146] buffer
x_and146 VSS VDD in[146] clk out[146] AND2x2_ASAP7_75t_SRAM
x_buf147 VDD VSS in[147] out[147] buffer
x_and147 VSS VDD in[147] clk out[147] AND2x2_ASAP7_75t_SRAM
x_buf148 VDD VSS in[148] out[148] buffer
x_and148 VSS VDD in[148] clk out[148] AND2x2_ASAP7_75t_SRAM
x_buf149 VDD VSS in[149] out[149] buffer
x_and149 VSS VDD in[149] clk out[149] AND2x2_ASAP7_75t_SRAM
x_buf150 VDD VSS in[150] out[150] buffer
x_and150 VSS VDD in[150] clk out[150] AND2x2_ASAP7_75t_SRAM
x_buf151 VDD VSS in[151] out[151] buffer
x_and151 VSS VDD in[151] clk out[151] AND2x2_ASAP7_75t_SRAM
x_buf152 VDD VSS in[152] out[152] buffer
x_and152 VSS VDD in[152] clk out[152] AND2x2_ASAP7_75t_SRAM
x_buf153 VDD VSS in[153] out[153] buffer
x_and153 VSS VDD in[153] clk out[153] AND2x2_ASAP7_75t_SRAM
x_buf154 VDD VSS in[154] out[154] buffer
x_and154 VSS VDD in[154] clk out[154] AND2x2_ASAP7_75t_SRAM
x_buf155 VDD VSS in[155] out[155] buffer
x_and155 VSS VDD in[155] clk out[155] AND2x2_ASAP7_75t_SRAM
x_buf156 VDD VSS in[156] out[156] buffer
x_and156 VSS VDD in[156] clk out[156] AND2x2_ASAP7_75t_SRAM
x_buf157 VDD VSS in[157] out[157] buffer
x_and157 VSS VDD in[157] clk out[157] AND2x2_ASAP7_75t_SRAM
x_buf158 VDD VSS in[158] out[158] buffer
x_and158 VSS VDD in[158] clk out[158] AND2x2_ASAP7_75t_SRAM
x_buf159 VDD VSS in[159] out[159] buffer
x_and159 VSS VDD in[159] clk out[159] AND2x2_ASAP7_75t_SRAM
x_buf160 VDD VSS in[160] out[160] buffer
x_and160 VSS VDD in[160] clk out[160] AND2x2_ASAP7_75t_SRAM
x_buf161 VDD VSS in[161] out[161] buffer
x_and161 VSS VDD in[161] clk out[161] AND2x2_ASAP7_75t_SRAM
x_buf162 VDD VSS in[162] out[162] buffer
x_and162 VSS VDD in[162] clk out[162] AND2x2_ASAP7_75t_SRAM
x_buf163 VDD VSS in[163] out[163] buffer
x_and163 VSS VDD in[163] clk out[163] AND2x2_ASAP7_75t_SRAM
x_buf164 VDD VSS in[164] out[164] buffer
x_and164 VSS VDD in[164] clk out[164] AND2x2_ASAP7_75t_SRAM
x_buf165 VDD VSS in[165] out[165] buffer
x_and165 VSS VDD in[165] clk out[165] AND2x2_ASAP7_75t_SRAM
x_buf166 VDD VSS in[166] out[166] buffer
x_and166 VSS VDD in[166] clk out[166] AND2x2_ASAP7_75t_SRAM
x_buf167 VDD VSS in[167] out[167] buffer
x_and167 VSS VDD in[167] clk out[167] AND2x2_ASAP7_75t_SRAM
x_buf168 VDD VSS in[168] out[168] buffer
x_and168 VSS VDD in[168] clk out[168] AND2x2_ASAP7_75t_SRAM
x_buf169 VDD VSS in[169] out[169] buffer
x_and169 VSS VDD in[169] clk out[169] AND2x2_ASAP7_75t_SRAM
x_buf170 VDD VSS in[170] out[170] buffer
x_and170 VSS VDD in[170] clk out[170] AND2x2_ASAP7_75t_SRAM
x_buf171 VDD VSS in[171] out[171] buffer
x_and171 VSS VDD in[171] clk out[171] AND2x2_ASAP7_75t_SRAM
x_buf172 VDD VSS in[172] out[172] buffer
x_and172 VSS VDD in[172] clk out[172] AND2x2_ASAP7_75t_SRAM
x_buf173 VDD VSS in[173] out[173] buffer
x_and173 VSS VDD in[173] clk out[173] AND2x2_ASAP7_75t_SRAM
x_buf174 VDD VSS in[174] out[174] buffer
x_and174 VSS VDD in[174] clk out[174] AND2x2_ASAP7_75t_SRAM
x_buf175 VDD VSS in[175] out[175] buffer
x_and175 VSS VDD in[175] clk out[175] AND2x2_ASAP7_75t_SRAM
x_buf176 VDD VSS in[176] out[176] buffer
x_and176 VSS VDD in[176] clk out[176] AND2x2_ASAP7_75t_SRAM
x_buf177 VDD VSS in[177] out[177] buffer
x_and177 VSS VDD in[177] clk out[177] AND2x2_ASAP7_75t_SRAM
x_buf178 VDD VSS in[178] out[178] buffer
x_and178 VSS VDD in[178] clk out[178] AND2x2_ASAP7_75t_SRAM
x_buf179 VDD VSS in[179] out[179] buffer
x_and179 VSS VDD in[179] clk out[179] AND2x2_ASAP7_75t_SRAM
x_buf180 VDD VSS in[180] out[180] buffer
x_and180 VSS VDD in[180] clk out[180] AND2x2_ASAP7_75t_SRAM
x_buf181 VDD VSS in[181] out[181] buffer
x_and181 VSS VDD in[181] clk out[181] AND2x2_ASAP7_75t_SRAM
x_buf182 VDD VSS in[182] out[182] buffer
x_and182 VSS VDD in[182] clk out[182] AND2x2_ASAP7_75t_SRAM
x_buf183 VDD VSS in[183] out[183] buffer
x_and183 VSS VDD in[183] clk out[183] AND2x2_ASAP7_75t_SRAM
x_buf184 VDD VSS in[184] out[184] buffer
x_and184 VSS VDD in[184] clk out[184] AND2x2_ASAP7_75t_SRAM
x_buf185 VDD VSS in[185] out[185] buffer
x_and185 VSS VDD in[185] clk out[185] AND2x2_ASAP7_75t_SRAM
x_buf186 VDD VSS in[186] out[186] buffer
x_and186 VSS VDD in[186] clk out[186] AND2x2_ASAP7_75t_SRAM
x_buf187 VDD VSS in[187] out[187] buffer
x_and187 VSS VDD in[187] clk out[187] AND2x2_ASAP7_75t_SRAM
x_buf188 VDD VSS in[188] out[188] buffer
x_and188 VSS VDD in[188] clk out[188] AND2x2_ASAP7_75t_SRAM
x_buf189 VDD VSS in[189] out[189] buffer
x_and189 VSS VDD in[189] clk out[189] AND2x2_ASAP7_75t_SRAM
x_buf190 VDD VSS in[190] out[190] buffer
x_and190 VSS VDD in[190] clk out[190] AND2x2_ASAP7_75t_SRAM
x_buf191 VDD VSS in[191] out[191] buffer
x_and191 VSS VDD in[191] clk out[191] AND2x2_ASAP7_75t_SRAM
x_buf192 VDD VSS in[192] out[192] buffer
x_and192 VSS VDD in[192] clk out[192] AND2x2_ASAP7_75t_SRAM
x_buf193 VDD VSS in[193] out[193] buffer
x_and193 VSS VDD in[193] clk out[193] AND2x2_ASAP7_75t_SRAM
x_buf194 VDD VSS in[194] out[194] buffer
x_and194 VSS VDD in[194] clk out[194] AND2x2_ASAP7_75t_SRAM
x_buf195 VDD VSS in[195] out[195] buffer
x_and195 VSS VDD in[195] clk out[195] AND2x2_ASAP7_75t_SRAM
x_buf196 VDD VSS in[196] out[196] buffer
x_and196 VSS VDD in[196] clk out[196] AND2x2_ASAP7_75t_SRAM
x_buf197 VDD VSS in[197] out[197] buffer
x_and197 VSS VDD in[197] clk out[197] AND2x2_ASAP7_75t_SRAM
x_buf198 VDD VSS in[198] out[198] buffer
x_and198 VSS VDD in[198] clk out[198] AND2x2_ASAP7_75t_SRAM
x_buf199 VDD VSS in[199] out[199] buffer
x_and199 VSS VDD in[199] clk out[199] AND2x2_ASAP7_75t_SRAM
x_buf200 VDD VSS in[200] out[200] buffer
x_and200 VSS VDD in[200] clk out[200] AND2x2_ASAP7_75t_SRAM
x_buf201 VDD VSS in[201] out[201] buffer
x_and201 VSS VDD in[201] clk out[201] AND2x2_ASAP7_75t_SRAM
x_buf202 VDD VSS in[202] out[202] buffer
x_and202 VSS VDD in[202] clk out[202] AND2x2_ASAP7_75t_SRAM
x_buf203 VDD VSS in[203] out[203] buffer
x_and203 VSS VDD in[203] clk out[203] AND2x2_ASAP7_75t_SRAM
x_buf204 VDD VSS in[204] out[204] buffer
x_and204 VSS VDD in[204] clk out[204] AND2x2_ASAP7_75t_SRAM
x_buf205 VDD VSS in[205] out[205] buffer
x_and205 VSS VDD in[205] clk out[205] AND2x2_ASAP7_75t_SRAM
x_buf206 VDD VSS in[206] out[206] buffer
x_and206 VSS VDD in[206] clk out[206] AND2x2_ASAP7_75t_SRAM
x_buf207 VDD VSS in[207] out[207] buffer
x_and207 VSS VDD in[207] clk out[207] AND2x2_ASAP7_75t_SRAM
x_buf208 VDD VSS in[208] out[208] buffer
x_and208 VSS VDD in[208] clk out[208] AND2x2_ASAP7_75t_SRAM
x_buf209 VDD VSS in[209] out[209] buffer
x_and209 VSS VDD in[209] clk out[209] AND2x2_ASAP7_75t_SRAM
x_buf210 VDD VSS in[210] out[210] buffer
x_and210 VSS VDD in[210] clk out[210] AND2x2_ASAP7_75t_SRAM
x_buf211 VDD VSS in[211] out[211] buffer
x_and211 VSS VDD in[211] clk out[211] AND2x2_ASAP7_75t_SRAM
x_buf212 VDD VSS in[212] out[212] buffer
x_and212 VSS VDD in[212] clk out[212] AND2x2_ASAP7_75t_SRAM
x_buf213 VDD VSS in[213] out[213] buffer
x_and213 VSS VDD in[213] clk out[213] AND2x2_ASAP7_75t_SRAM
x_buf214 VDD VSS in[214] out[214] buffer
x_and214 VSS VDD in[214] clk out[214] AND2x2_ASAP7_75t_SRAM
x_buf215 VDD VSS in[215] out[215] buffer
x_and215 VSS VDD in[215] clk out[215] AND2x2_ASAP7_75t_SRAM
x_buf216 VDD VSS in[216] out[216] buffer
x_and216 VSS VDD in[216] clk out[216] AND2x2_ASAP7_75t_SRAM
x_buf217 VDD VSS in[217] out[217] buffer
x_and217 VSS VDD in[217] clk out[217] AND2x2_ASAP7_75t_SRAM
x_buf218 VDD VSS in[218] out[218] buffer
x_and218 VSS VDD in[218] clk out[218] AND2x2_ASAP7_75t_SRAM
x_buf219 VDD VSS in[219] out[219] buffer
x_and219 VSS VDD in[219] clk out[219] AND2x2_ASAP7_75t_SRAM
x_buf220 VDD VSS in[220] out[220] buffer
x_and220 VSS VDD in[220] clk out[220] AND2x2_ASAP7_75t_SRAM
x_buf221 VDD VSS in[221] out[221] buffer
x_and221 VSS VDD in[221] clk out[221] AND2x2_ASAP7_75t_SRAM
x_buf222 VDD VSS in[222] out[222] buffer
x_and222 VSS VDD in[222] clk out[222] AND2x2_ASAP7_75t_SRAM
x_buf223 VDD VSS in[223] out[223] buffer
x_and223 VSS VDD in[223] clk out[223] AND2x2_ASAP7_75t_SRAM
x_buf224 VDD VSS in[224] out[224] buffer
x_and224 VSS VDD in[224] clk out[224] AND2x2_ASAP7_75t_SRAM
x_buf225 VDD VSS in[225] out[225] buffer
x_and225 VSS VDD in[225] clk out[225] AND2x2_ASAP7_75t_SRAM
x_buf226 VDD VSS in[226] out[226] buffer
x_and226 VSS VDD in[226] clk out[226] AND2x2_ASAP7_75t_SRAM
x_buf227 VDD VSS in[227] out[227] buffer
x_and227 VSS VDD in[227] clk out[227] AND2x2_ASAP7_75t_SRAM
x_buf228 VDD VSS in[228] out[228] buffer
x_and228 VSS VDD in[228] clk out[228] AND2x2_ASAP7_75t_SRAM
x_buf229 VDD VSS in[229] out[229] buffer
x_and229 VSS VDD in[229] clk out[229] AND2x2_ASAP7_75t_SRAM
x_buf230 VDD VSS in[230] out[230] buffer
x_and230 VSS VDD in[230] clk out[230] AND2x2_ASAP7_75t_SRAM
x_buf231 VDD VSS in[231] out[231] buffer
x_and231 VSS VDD in[231] clk out[231] AND2x2_ASAP7_75t_SRAM
x_buf232 VDD VSS in[232] out[232] buffer
x_and232 VSS VDD in[232] clk out[232] AND2x2_ASAP7_75t_SRAM
x_buf233 VDD VSS in[233] out[233] buffer
x_and233 VSS VDD in[233] clk out[233] AND2x2_ASAP7_75t_SRAM
x_buf234 VDD VSS in[234] out[234] buffer
x_and234 VSS VDD in[234] clk out[234] AND2x2_ASAP7_75t_SRAM
x_buf235 VDD VSS in[235] out[235] buffer
x_and235 VSS VDD in[235] clk out[235] AND2x2_ASAP7_75t_SRAM
x_buf236 VDD VSS in[236] out[236] buffer
x_and236 VSS VDD in[236] clk out[236] AND2x2_ASAP7_75t_SRAM
x_buf237 VDD VSS in[237] out[237] buffer
x_and237 VSS VDD in[237] clk out[237] AND2x2_ASAP7_75t_SRAM
x_buf238 VDD VSS in[238] out[238] buffer
x_and238 VSS VDD in[238] clk out[238] AND2x2_ASAP7_75t_SRAM
x_buf239 VDD VSS in[239] out[239] buffer
x_and239 VSS VDD in[239] clk out[239] AND2x2_ASAP7_75t_SRAM
x_buf240 VDD VSS in[240] out[240] buffer
x_and240 VSS VDD in[240] clk out[240] AND2x2_ASAP7_75t_SRAM
x_buf241 VDD VSS in[241] out[241] buffer
x_and241 VSS VDD in[241] clk out[241] AND2x2_ASAP7_75t_SRAM
x_buf242 VDD VSS in[242] out[242] buffer
x_and242 VSS VDD in[242] clk out[242] AND2x2_ASAP7_75t_SRAM
x_buf243 VDD VSS in[243] out[243] buffer
x_and243 VSS VDD in[243] clk out[243] AND2x2_ASAP7_75t_SRAM
x_buf244 VDD VSS in[244] out[244] buffer
x_and244 VSS VDD in[244] clk out[244] AND2x2_ASAP7_75t_SRAM
x_buf245 VDD VSS in[245] out[245] buffer
x_and245 VSS VDD in[245] clk out[245] AND2x2_ASAP7_75t_SRAM
x_buf246 VDD VSS in[246] out[246] buffer
x_and246 VSS VDD in[246] clk out[246] AND2x2_ASAP7_75t_SRAM
x_buf247 VDD VSS in[247] out[247] buffer
x_and247 VSS VDD in[247] clk out[247] AND2x2_ASAP7_75t_SRAM
x_buf248 VDD VSS in[248] out[248] buffer
x_and248 VSS VDD in[248] clk out[248] AND2x2_ASAP7_75t_SRAM
x_buf249 VDD VSS in[249] out[249] buffer
x_and249 VSS VDD in[249] clk out[249] AND2x2_ASAP7_75t_SRAM
x_buf250 VDD VSS in[250] out[250] buffer
x_and250 VSS VDD in[250] clk out[250] AND2x2_ASAP7_75t_SRAM
x_buf251 VDD VSS in[251] out[251] buffer
x_and251 VSS VDD in[251] clk out[251] AND2x2_ASAP7_75t_SRAM
x_buf252 VDD VSS in[252] out[252] buffer
x_and252 VSS VDD in[252] clk out[252] AND2x2_ASAP7_75t_SRAM
x_buf253 VDD VSS in[253] out[253] buffer
x_and253 VSS VDD in[253] clk out[253] AND2x2_ASAP7_75t_SRAM
x_buf254 VDD VSS in[254] out[254] buffer
x_and254 VSS VDD in[254] clk out[254] AND2x2_ASAP7_75t_SRAM
x_buf255 VDD VSS in[255] out[255] buffer
x_and255 VSS VDD in[255] clk out[255] AND2x2_ASAP7_75t_SRAM
x_buf256 VDD VSS in[256] out[256] buffer
x_and256 VSS VDD in[256] clk out[256] AND2x2_ASAP7_75t_SRAM
x_buf257 VDD VSS in[257] out[257] buffer
x_and257 VSS VDD in[257] clk out[257] AND2x2_ASAP7_75t_SRAM
x_buf258 VDD VSS in[258] out[258] buffer
x_and258 VSS VDD in[258] clk out[258] AND2x2_ASAP7_75t_SRAM
x_buf259 VDD VSS in[259] out[259] buffer
x_and259 VSS VDD in[259] clk out[259] AND2x2_ASAP7_75t_SRAM
x_buf260 VDD VSS in[260] out[260] buffer
x_and260 VSS VDD in[260] clk out[260] AND2x2_ASAP7_75t_SRAM
x_buf261 VDD VSS in[261] out[261] buffer
x_and261 VSS VDD in[261] clk out[261] AND2x2_ASAP7_75t_SRAM
x_buf262 VDD VSS in[262] out[262] buffer
x_and262 VSS VDD in[262] clk out[262] AND2x2_ASAP7_75t_SRAM
x_buf263 VDD VSS in[263] out[263] buffer
x_and263 VSS VDD in[263] clk out[263] AND2x2_ASAP7_75t_SRAM
x_buf264 VDD VSS in[264] out[264] buffer
x_and264 VSS VDD in[264] clk out[264] AND2x2_ASAP7_75t_SRAM
x_buf265 VDD VSS in[265] out[265] buffer
x_and265 VSS VDD in[265] clk out[265] AND2x2_ASAP7_75t_SRAM
x_buf266 VDD VSS in[266] out[266] buffer
x_and266 VSS VDD in[266] clk out[266] AND2x2_ASAP7_75t_SRAM
x_buf267 VDD VSS in[267] out[267] buffer
x_and267 VSS VDD in[267] clk out[267] AND2x2_ASAP7_75t_SRAM
x_buf268 VDD VSS in[268] out[268] buffer
x_and268 VSS VDD in[268] clk out[268] AND2x2_ASAP7_75t_SRAM
x_buf269 VDD VSS in[269] out[269] buffer
x_and269 VSS VDD in[269] clk out[269] AND2x2_ASAP7_75t_SRAM
x_buf270 VDD VSS in[270] out[270] buffer
x_and270 VSS VDD in[270] clk out[270] AND2x2_ASAP7_75t_SRAM
x_buf271 VDD VSS in[271] out[271] buffer
x_and271 VSS VDD in[271] clk out[271] AND2x2_ASAP7_75t_SRAM
x_buf272 VDD VSS in[272] out[272] buffer
x_and272 VSS VDD in[272] clk out[272] AND2x2_ASAP7_75t_SRAM
x_buf273 VDD VSS in[273] out[273] buffer
x_and273 VSS VDD in[273] clk out[273] AND2x2_ASAP7_75t_SRAM
x_buf274 VDD VSS in[274] out[274] buffer
x_and274 VSS VDD in[274] clk out[274] AND2x2_ASAP7_75t_SRAM
x_buf275 VDD VSS in[275] out[275] buffer
x_and275 VSS VDD in[275] clk out[275] AND2x2_ASAP7_75t_SRAM
x_buf276 VDD VSS in[276] out[276] buffer
x_and276 VSS VDD in[276] clk out[276] AND2x2_ASAP7_75t_SRAM
x_buf277 VDD VSS in[277] out[277] buffer
x_and277 VSS VDD in[277] clk out[277] AND2x2_ASAP7_75t_SRAM
x_buf278 VDD VSS in[278] out[278] buffer
x_and278 VSS VDD in[278] clk out[278] AND2x2_ASAP7_75t_SRAM
x_buf279 VDD VSS in[279] out[279] buffer
x_and279 VSS VDD in[279] clk out[279] AND2x2_ASAP7_75t_SRAM
x_buf280 VDD VSS in[280] out[280] buffer
x_and280 VSS VDD in[280] clk out[280] AND2x2_ASAP7_75t_SRAM
x_buf281 VDD VSS in[281] out[281] buffer
x_and281 VSS VDD in[281] clk out[281] AND2x2_ASAP7_75t_SRAM
x_buf282 VDD VSS in[282] out[282] buffer
x_and282 VSS VDD in[282] clk out[282] AND2x2_ASAP7_75t_SRAM
x_buf283 VDD VSS in[283] out[283] buffer
x_and283 VSS VDD in[283] clk out[283] AND2x2_ASAP7_75t_SRAM
x_buf284 VDD VSS in[284] out[284] buffer
x_and284 VSS VDD in[284] clk out[284] AND2x2_ASAP7_75t_SRAM
x_buf285 VDD VSS in[285] out[285] buffer
x_and285 VSS VDD in[285] clk out[285] AND2x2_ASAP7_75t_SRAM
x_buf286 VDD VSS in[286] out[286] buffer
x_and286 VSS VDD in[286] clk out[286] AND2x2_ASAP7_75t_SRAM
x_buf287 VDD VSS in[287] out[287] buffer
x_and287 VSS VDD in[287] clk out[287] AND2x2_ASAP7_75t_SRAM
x_buf288 VDD VSS in[288] out[288] buffer
x_and288 VSS VDD in[288] clk out[288] AND2x2_ASAP7_75t_SRAM
x_buf289 VDD VSS in[289] out[289] buffer
x_and289 VSS VDD in[289] clk out[289] AND2x2_ASAP7_75t_SRAM
x_buf290 VDD VSS in[290] out[290] buffer
x_and290 VSS VDD in[290] clk out[290] AND2x2_ASAP7_75t_SRAM
x_buf291 VDD VSS in[291] out[291] buffer
x_and291 VSS VDD in[291] clk out[291] AND2x2_ASAP7_75t_SRAM
x_buf292 VDD VSS in[292] out[292] buffer
x_and292 VSS VDD in[292] clk out[292] AND2x2_ASAP7_75t_SRAM
x_buf293 VDD VSS in[293] out[293] buffer
x_and293 VSS VDD in[293] clk out[293] AND2x2_ASAP7_75t_SRAM
x_buf294 VDD VSS in[294] out[294] buffer
x_and294 VSS VDD in[294] clk out[294] AND2x2_ASAP7_75t_SRAM
x_buf295 VDD VSS in[295] out[295] buffer
x_and295 VSS VDD in[295] clk out[295] AND2x2_ASAP7_75t_SRAM
x_buf296 VDD VSS in[296] out[296] buffer
x_and296 VSS VDD in[296] clk out[296] AND2x2_ASAP7_75t_SRAM
x_buf297 VDD VSS in[297] out[297] buffer
x_and297 VSS VDD in[297] clk out[297] AND2x2_ASAP7_75t_SRAM
x_buf298 VDD VSS in[298] out[298] buffer
x_and298 VSS VDD in[298] clk out[298] AND2x2_ASAP7_75t_SRAM
x_buf299 VDD VSS in[299] out[299] buffer
x_and299 VSS VDD in[299] clk out[299] AND2x2_ASAP7_75t_SRAM
x_buf300 VDD VSS in[300] out[300] buffer
x_and300 VSS VDD in[300] clk out[300] AND2x2_ASAP7_75t_SRAM
x_buf301 VDD VSS in[301] out[301] buffer
x_and301 VSS VDD in[301] clk out[301] AND2x2_ASAP7_75t_SRAM
x_buf302 VDD VSS in[302] out[302] buffer
x_and302 VSS VDD in[302] clk out[302] AND2x2_ASAP7_75t_SRAM
x_buf303 VDD VSS in[303] out[303] buffer
x_and303 VSS VDD in[303] clk out[303] AND2x2_ASAP7_75t_SRAM
x_buf304 VDD VSS in[304] out[304] buffer
x_and304 VSS VDD in[304] clk out[304] AND2x2_ASAP7_75t_SRAM
x_buf305 VDD VSS in[305] out[305] buffer
x_and305 VSS VDD in[305] clk out[305] AND2x2_ASAP7_75t_SRAM
x_buf306 VDD VSS in[306] out[306] buffer
x_and306 VSS VDD in[306] clk out[306] AND2x2_ASAP7_75t_SRAM
x_buf307 VDD VSS in[307] out[307] buffer
x_and307 VSS VDD in[307] clk out[307] AND2x2_ASAP7_75t_SRAM
x_buf308 VDD VSS in[308] out[308] buffer
x_and308 VSS VDD in[308] clk out[308] AND2x2_ASAP7_75t_SRAM
x_buf309 VDD VSS in[309] out[309] buffer
x_and309 VSS VDD in[309] clk out[309] AND2x2_ASAP7_75t_SRAM
x_buf310 VDD VSS in[310] out[310] buffer
x_and310 VSS VDD in[310] clk out[310] AND2x2_ASAP7_75t_SRAM
x_buf311 VDD VSS in[311] out[311] buffer
x_and311 VSS VDD in[311] clk out[311] AND2x2_ASAP7_75t_SRAM
x_buf312 VDD VSS in[312] out[312] buffer
x_and312 VSS VDD in[312] clk out[312] AND2x2_ASAP7_75t_SRAM
x_buf313 VDD VSS in[313] out[313] buffer
x_and313 VSS VDD in[313] clk out[313] AND2x2_ASAP7_75t_SRAM
x_buf314 VDD VSS in[314] out[314] buffer
x_and314 VSS VDD in[314] clk out[314] AND2x2_ASAP7_75t_SRAM
x_buf315 VDD VSS in[315] out[315] buffer
x_and315 VSS VDD in[315] clk out[315] AND2x2_ASAP7_75t_SRAM
x_buf316 VDD VSS in[316] out[316] buffer
x_and316 VSS VDD in[316] clk out[316] AND2x2_ASAP7_75t_SRAM
x_buf317 VDD VSS in[317] out[317] buffer
x_and317 VSS VDD in[317] clk out[317] AND2x2_ASAP7_75t_SRAM
x_buf318 VDD VSS in[318] out[318] buffer
x_and318 VSS VDD in[318] clk out[318] AND2x2_ASAP7_75t_SRAM
x_buf319 VDD VSS in[319] out[319] buffer
x_and319 VSS VDD in[319] clk out[319] AND2x2_ASAP7_75t_SRAM
x_buf320 VDD VSS in[320] out[320] buffer
x_and320 VSS VDD in[320] clk out[320] AND2x2_ASAP7_75t_SRAM
x_buf321 VDD VSS in[321] out[321] buffer
x_and321 VSS VDD in[321] clk out[321] AND2x2_ASAP7_75t_SRAM
x_buf322 VDD VSS in[322] out[322] buffer
x_and322 VSS VDD in[322] clk out[322] AND2x2_ASAP7_75t_SRAM
x_buf323 VDD VSS in[323] out[323] buffer
x_and323 VSS VDD in[323] clk out[323] AND2x2_ASAP7_75t_SRAM
x_buf324 VDD VSS in[324] out[324] buffer
x_and324 VSS VDD in[324] clk out[324] AND2x2_ASAP7_75t_SRAM
x_buf325 VDD VSS in[325] out[325] buffer
x_and325 VSS VDD in[325] clk out[325] AND2x2_ASAP7_75t_SRAM
x_buf326 VDD VSS in[326] out[326] buffer
x_and326 VSS VDD in[326] clk out[326] AND2x2_ASAP7_75t_SRAM
x_buf327 VDD VSS in[327] out[327] buffer
x_and327 VSS VDD in[327] clk out[327] AND2x2_ASAP7_75t_SRAM
x_buf328 VDD VSS in[328] out[328] buffer
x_and328 VSS VDD in[328] clk out[328] AND2x2_ASAP7_75t_SRAM
x_buf329 VDD VSS in[329] out[329] buffer
x_and329 VSS VDD in[329] clk out[329] AND2x2_ASAP7_75t_SRAM
x_buf330 VDD VSS in[330] out[330] buffer
x_and330 VSS VDD in[330] clk out[330] AND2x2_ASAP7_75t_SRAM
x_buf331 VDD VSS in[331] out[331] buffer
x_and331 VSS VDD in[331] clk out[331] AND2x2_ASAP7_75t_SRAM
x_buf332 VDD VSS in[332] out[332] buffer
x_and332 VSS VDD in[332] clk out[332] AND2x2_ASAP7_75t_SRAM
x_buf333 VDD VSS in[333] out[333] buffer
x_and333 VSS VDD in[333] clk out[333] AND2x2_ASAP7_75t_SRAM
x_buf334 VDD VSS in[334] out[334] buffer
x_and334 VSS VDD in[334] clk out[334] AND2x2_ASAP7_75t_SRAM
x_buf335 VDD VSS in[335] out[335] buffer
x_and335 VSS VDD in[335] clk out[335] AND2x2_ASAP7_75t_SRAM
x_buf336 VDD VSS in[336] out[336] buffer
x_and336 VSS VDD in[336] clk out[336] AND2x2_ASAP7_75t_SRAM
x_buf337 VDD VSS in[337] out[337] buffer
x_and337 VSS VDD in[337] clk out[337] AND2x2_ASAP7_75t_SRAM
x_buf338 VDD VSS in[338] out[338] buffer
x_and338 VSS VDD in[338] clk out[338] AND2x2_ASAP7_75t_SRAM
x_buf339 VDD VSS in[339] out[339] buffer
x_and339 VSS VDD in[339] clk out[339] AND2x2_ASAP7_75t_SRAM
x_buf340 VDD VSS in[340] out[340] buffer
x_and340 VSS VDD in[340] clk out[340] AND2x2_ASAP7_75t_SRAM
x_buf341 VDD VSS in[341] out[341] buffer
x_and341 VSS VDD in[341] clk out[341] AND2x2_ASAP7_75t_SRAM
x_buf342 VDD VSS in[342] out[342] buffer
x_and342 VSS VDD in[342] clk out[342] AND2x2_ASAP7_75t_SRAM
x_buf343 VDD VSS in[343] out[343] buffer
x_and343 VSS VDD in[343] clk out[343] AND2x2_ASAP7_75t_SRAM
x_buf344 VDD VSS in[344] out[344] buffer
x_and344 VSS VDD in[344] clk out[344] AND2x2_ASAP7_75t_SRAM
x_buf345 VDD VSS in[345] out[345] buffer
x_and345 VSS VDD in[345] clk out[345] AND2x2_ASAP7_75t_SRAM
x_buf346 VDD VSS in[346] out[346] buffer
x_and346 VSS VDD in[346] clk out[346] AND2x2_ASAP7_75t_SRAM
x_buf347 VDD VSS in[347] out[347] buffer
x_and347 VSS VDD in[347] clk out[347] AND2x2_ASAP7_75t_SRAM
x_buf348 VDD VSS in[348] out[348] buffer
x_and348 VSS VDD in[348] clk out[348] AND2x2_ASAP7_75t_SRAM
x_buf349 VDD VSS in[349] out[349] buffer
x_and349 VSS VDD in[349] clk out[349] AND2x2_ASAP7_75t_SRAM
x_buf350 VDD VSS in[350] out[350] buffer
x_and350 VSS VDD in[350] clk out[350] AND2x2_ASAP7_75t_SRAM
x_buf351 VDD VSS in[351] out[351] buffer
x_and351 VSS VDD in[351] clk out[351] AND2x2_ASAP7_75t_SRAM
x_buf352 VDD VSS in[352] out[352] buffer
x_and352 VSS VDD in[352] clk out[352] AND2x2_ASAP7_75t_SRAM
x_buf353 VDD VSS in[353] out[353] buffer
x_and353 VSS VDD in[353] clk out[353] AND2x2_ASAP7_75t_SRAM
x_buf354 VDD VSS in[354] out[354] buffer
x_and354 VSS VDD in[354] clk out[354] AND2x2_ASAP7_75t_SRAM
x_buf355 VDD VSS in[355] out[355] buffer
x_and355 VSS VDD in[355] clk out[355] AND2x2_ASAP7_75t_SRAM
x_buf356 VDD VSS in[356] out[356] buffer
x_and356 VSS VDD in[356] clk out[356] AND2x2_ASAP7_75t_SRAM
x_buf357 VDD VSS in[357] out[357] buffer
x_and357 VSS VDD in[357] clk out[357] AND2x2_ASAP7_75t_SRAM
x_buf358 VDD VSS in[358] out[358] buffer
x_and358 VSS VDD in[358] clk out[358] AND2x2_ASAP7_75t_SRAM
x_buf359 VDD VSS in[359] out[359] buffer
x_and359 VSS VDD in[359] clk out[359] AND2x2_ASAP7_75t_SRAM
x_buf360 VDD VSS in[360] out[360] buffer
x_and360 VSS VDD in[360] clk out[360] AND2x2_ASAP7_75t_SRAM
x_buf361 VDD VSS in[361] out[361] buffer
x_and361 VSS VDD in[361] clk out[361] AND2x2_ASAP7_75t_SRAM
x_buf362 VDD VSS in[362] out[362] buffer
x_and362 VSS VDD in[362] clk out[362] AND2x2_ASAP7_75t_SRAM
x_buf363 VDD VSS in[363] out[363] buffer
x_and363 VSS VDD in[363] clk out[363] AND2x2_ASAP7_75t_SRAM
x_buf364 VDD VSS in[364] out[364] buffer
x_and364 VSS VDD in[364] clk out[364] AND2x2_ASAP7_75t_SRAM
x_buf365 VDD VSS in[365] out[365] buffer
x_and365 VSS VDD in[365] clk out[365] AND2x2_ASAP7_75t_SRAM
x_buf366 VDD VSS in[366] out[366] buffer
x_and366 VSS VDD in[366] clk out[366] AND2x2_ASAP7_75t_SRAM
x_buf367 VDD VSS in[367] out[367] buffer
x_and367 VSS VDD in[367] clk out[367] AND2x2_ASAP7_75t_SRAM
x_buf368 VDD VSS in[368] out[368] buffer
x_and368 VSS VDD in[368] clk out[368] AND2x2_ASAP7_75t_SRAM
x_buf369 VDD VSS in[369] out[369] buffer
x_and369 VSS VDD in[369] clk out[369] AND2x2_ASAP7_75t_SRAM
x_buf370 VDD VSS in[370] out[370] buffer
x_and370 VSS VDD in[370] clk out[370] AND2x2_ASAP7_75t_SRAM
x_buf371 VDD VSS in[371] out[371] buffer
x_and371 VSS VDD in[371] clk out[371] AND2x2_ASAP7_75t_SRAM
x_buf372 VDD VSS in[372] out[372] buffer
x_and372 VSS VDD in[372] clk out[372] AND2x2_ASAP7_75t_SRAM
x_buf373 VDD VSS in[373] out[373] buffer
x_and373 VSS VDD in[373] clk out[373] AND2x2_ASAP7_75t_SRAM
x_buf374 VDD VSS in[374] out[374] buffer
x_and374 VSS VDD in[374] clk out[374] AND2x2_ASAP7_75t_SRAM
x_buf375 VDD VSS in[375] out[375] buffer
x_and375 VSS VDD in[375] clk out[375] AND2x2_ASAP7_75t_SRAM
x_buf376 VDD VSS in[376] out[376] buffer
x_and376 VSS VDD in[376] clk out[376] AND2x2_ASAP7_75t_SRAM
x_buf377 VDD VSS in[377] out[377] buffer
x_and377 VSS VDD in[377] clk out[377] AND2x2_ASAP7_75t_SRAM
x_buf378 VDD VSS in[378] out[378] buffer
x_and378 VSS VDD in[378] clk out[378] AND2x2_ASAP7_75t_SRAM
x_buf379 VDD VSS in[379] out[379] buffer
x_and379 VSS VDD in[379] clk out[379] AND2x2_ASAP7_75t_SRAM
x_buf380 VDD VSS in[380] out[380] buffer
x_and380 VSS VDD in[380] clk out[380] AND2x2_ASAP7_75t_SRAM
x_buf381 VDD VSS in[381] out[381] buffer
x_and381 VSS VDD in[381] clk out[381] AND2x2_ASAP7_75t_SRAM
x_buf382 VDD VSS in[382] out[382] buffer
x_and382 VSS VDD in[382] clk out[382] AND2x2_ASAP7_75t_SRAM
x_buf383 VDD VSS in[383] out[383] buffer
x_and383 VSS VDD in[383] clk out[383] AND2x2_ASAP7_75t_SRAM
x_buf384 VDD VSS in[384] out[384] buffer
x_and384 VSS VDD in[384] clk out[384] AND2x2_ASAP7_75t_SRAM
x_buf385 VDD VSS in[385] out[385] buffer
x_and385 VSS VDD in[385] clk out[385] AND2x2_ASAP7_75t_SRAM
x_buf386 VDD VSS in[386] out[386] buffer
x_and386 VSS VDD in[386] clk out[386] AND2x2_ASAP7_75t_SRAM
x_buf387 VDD VSS in[387] out[387] buffer
x_and387 VSS VDD in[387] clk out[387] AND2x2_ASAP7_75t_SRAM
x_buf388 VDD VSS in[388] out[388] buffer
x_and388 VSS VDD in[388] clk out[388] AND2x2_ASAP7_75t_SRAM
x_buf389 VDD VSS in[389] out[389] buffer
x_and389 VSS VDD in[389] clk out[389] AND2x2_ASAP7_75t_SRAM
x_buf390 VDD VSS in[390] out[390] buffer
x_and390 VSS VDD in[390] clk out[390] AND2x2_ASAP7_75t_SRAM
x_buf391 VDD VSS in[391] out[391] buffer
x_and391 VSS VDD in[391] clk out[391] AND2x2_ASAP7_75t_SRAM
x_buf392 VDD VSS in[392] out[392] buffer
x_and392 VSS VDD in[392] clk out[392] AND2x2_ASAP7_75t_SRAM
x_buf393 VDD VSS in[393] out[393] buffer
x_and393 VSS VDD in[393] clk out[393] AND2x2_ASAP7_75t_SRAM
x_buf394 VDD VSS in[394] out[394] buffer
x_and394 VSS VDD in[394] clk out[394] AND2x2_ASAP7_75t_SRAM
x_buf395 VDD VSS in[395] out[395] buffer
x_and395 VSS VDD in[395] clk out[395] AND2x2_ASAP7_75t_SRAM
x_buf396 VDD VSS in[396] out[396] buffer
x_and396 VSS VDD in[396] clk out[396] AND2x2_ASAP7_75t_SRAM
x_buf397 VDD VSS in[397] out[397] buffer
x_and397 VSS VDD in[397] clk out[397] AND2x2_ASAP7_75t_SRAM
x_buf398 VDD VSS in[398] out[398] buffer
x_and398 VSS VDD in[398] clk out[398] AND2x2_ASAP7_75t_SRAM
x_buf399 VDD VSS in[399] out[399] buffer
x_and399 VSS VDD in[399] clk out[399] AND2x2_ASAP7_75t_SRAM
x_buf400 VDD VSS in[400] out[400] buffer
x_and400 VSS VDD in[400] clk out[400] AND2x2_ASAP7_75t_SRAM
x_buf401 VDD VSS in[401] out[401] buffer
x_and401 VSS VDD in[401] clk out[401] AND2x2_ASAP7_75t_SRAM
x_buf402 VDD VSS in[402] out[402] buffer
x_and402 VSS VDD in[402] clk out[402] AND2x2_ASAP7_75t_SRAM
x_buf403 VDD VSS in[403] out[403] buffer
x_and403 VSS VDD in[403] clk out[403] AND2x2_ASAP7_75t_SRAM
x_buf404 VDD VSS in[404] out[404] buffer
x_and404 VSS VDD in[404] clk out[404] AND2x2_ASAP7_75t_SRAM
x_buf405 VDD VSS in[405] out[405] buffer
x_and405 VSS VDD in[405] clk out[405] AND2x2_ASAP7_75t_SRAM
x_buf406 VDD VSS in[406] out[406] buffer
x_and406 VSS VDD in[406] clk out[406] AND2x2_ASAP7_75t_SRAM
x_buf407 VDD VSS in[407] out[407] buffer
x_and407 VSS VDD in[407] clk out[407] AND2x2_ASAP7_75t_SRAM
x_buf408 VDD VSS in[408] out[408] buffer
x_and408 VSS VDD in[408] clk out[408] AND2x2_ASAP7_75t_SRAM
x_buf409 VDD VSS in[409] out[409] buffer
x_and409 VSS VDD in[409] clk out[409] AND2x2_ASAP7_75t_SRAM
x_buf410 VDD VSS in[410] out[410] buffer
x_and410 VSS VDD in[410] clk out[410] AND2x2_ASAP7_75t_SRAM
x_buf411 VDD VSS in[411] out[411] buffer
x_and411 VSS VDD in[411] clk out[411] AND2x2_ASAP7_75t_SRAM
x_buf412 VDD VSS in[412] out[412] buffer
x_and412 VSS VDD in[412] clk out[412] AND2x2_ASAP7_75t_SRAM
x_buf413 VDD VSS in[413] out[413] buffer
x_and413 VSS VDD in[413] clk out[413] AND2x2_ASAP7_75t_SRAM
x_buf414 VDD VSS in[414] out[414] buffer
x_and414 VSS VDD in[414] clk out[414] AND2x2_ASAP7_75t_SRAM
x_buf415 VDD VSS in[415] out[415] buffer
x_and415 VSS VDD in[415] clk out[415] AND2x2_ASAP7_75t_SRAM
x_buf416 VDD VSS in[416] out[416] buffer
x_and416 VSS VDD in[416] clk out[416] AND2x2_ASAP7_75t_SRAM
x_buf417 VDD VSS in[417] out[417] buffer
x_and417 VSS VDD in[417] clk out[417] AND2x2_ASAP7_75t_SRAM
x_buf418 VDD VSS in[418] out[418] buffer
x_and418 VSS VDD in[418] clk out[418] AND2x2_ASAP7_75t_SRAM
x_buf419 VDD VSS in[419] out[419] buffer
x_and419 VSS VDD in[419] clk out[419] AND2x2_ASAP7_75t_SRAM
x_buf420 VDD VSS in[420] out[420] buffer
x_and420 VSS VDD in[420] clk out[420] AND2x2_ASAP7_75t_SRAM
x_buf421 VDD VSS in[421] out[421] buffer
x_and421 VSS VDD in[421] clk out[421] AND2x2_ASAP7_75t_SRAM
x_buf422 VDD VSS in[422] out[422] buffer
x_and422 VSS VDD in[422] clk out[422] AND2x2_ASAP7_75t_SRAM
x_buf423 VDD VSS in[423] out[423] buffer
x_and423 VSS VDD in[423] clk out[423] AND2x2_ASAP7_75t_SRAM
x_buf424 VDD VSS in[424] out[424] buffer
x_and424 VSS VDD in[424] clk out[424] AND2x2_ASAP7_75t_SRAM
x_buf425 VDD VSS in[425] out[425] buffer
x_and425 VSS VDD in[425] clk out[425] AND2x2_ASAP7_75t_SRAM
x_buf426 VDD VSS in[426] out[426] buffer
x_and426 VSS VDD in[426] clk out[426] AND2x2_ASAP7_75t_SRAM
x_buf427 VDD VSS in[427] out[427] buffer
x_and427 VSS VDD in[427] clk out[427] AND2x2_ASAP7_75t_SRAM
x_buf428 VDD VSS in[428] out[428] buffer
x_and428 VSS VDD in[428] clk out[428] AND2x2_ASAP7_75t_SRAM
x_buf429 VDD VSS in[429] out[429] buffer
x_and429 VSS VDD in[429] clk out[429] AND2x2_ASAP7_75t_SRAM
x_buf430 VDD VSS in[430] out[430] buffer
x_and430 VSS VDD in[430] clk out[430] AND2x2_ASAP7_75t_SRAM
x_buf431 VDD VSS in[431] out[431] buffer
x_and431 VSS VDD in[431] clk out[431] AND2x2_ASAP7_75t_SRAM
x_buf432 VDD VSS in[432] out[432] buffer
x_and432 VSS VDD in[432] clk out[432] AND2x2_ASAP7_75t_SRAM
x_buf433 VDD VSS in[433] out[433] buffer
x_and433 VSS VDD in[433] clk out[433] AND2x2_ASAP7_75t_SRAM
x_buf434 VDD VSS in[434] out[434] buffer
x_and434 VSS VDD in[434] clk out[434] AND2x2_ASAP7_75t_SRAM
x_buf435 VDD VSS in[435] out[435] buffer
x_and435 VSS VDD in[435] clk out[435] AND2x2_ASAP7_75t_SRAM
x_buf436 VDD VSS in[436] out[436] buffer
x_and436 VSS VDD in[436] clk out[436] AND2x2_ASAP7_75t_SRAM
x_buf437 VDD VSS in[437] out[437] buffer
x_and437 VSS VDD in[437] clk out[437] AND2x2_ASAP7_75t_SRAM
x_buf438 VDD VSS in[438] out[438] buffer
x_and438 VSS VDD in[438] clk out[438] AND2x2_ASAP7_75t_SRAM
x_buf439 VDD VSS in[439] out[439] buffer
x_and439 VSS VDD in[439] clk out[439] AND2x2_ASAP7_75t_SRAM
x_buf440 VDD VSS in[440] out[440] buffer
x_and440 VSS VDD in[440] clk out[440] AND2x2_ASAP7_75t_SRAM
x_buf441 VDD VSS in[441] out[441] buffer
x_and441 VSS VDD in[441] clk out[441] AND2x2_ASAP7_75t_SRAM
x_buf442 VDD VSS in[442] out[442] buffer
x_and442 VSS VDD in[442] clk out[442] AND2x2_ASAP7_75t_SRAM
x_buf443 VDD VSS in[443] out[443] buffer
x_and443 VSS VDD in[443] clk out[443] AND2x2_ASAP7_75t_SRAM
x_buf444 VDD VSS in[444] out[444] buffer
x_and444 VSS VDD in[444] clk out[444] AND2x2_ASAP7_75t_SRAM
x_buf445 VDD VSS in[445] out[445] buffer
x_and445 VSS VDD in[445] clk out[445] AND2x2_ASAP7_75t_SRAM
x_buf446 VDD VSS in[446] out[446] buffer
x_and446 VSS VDD in[446] clk out[446] AND2x2_ASAP7_75t_SRAM
x_buf447 VDD VSS in[447] out[447] buffer
x_and447 VSS VDD in[447] clk out[447] AND2x2_ASAP7_75t_SRAM
x_buf448 VDD VSS in[448] out[448] buffer
x_and448 VSS VDD in[448] clk out[448] AND2x2_ASAP7_75t_SRAM
x_buf449 VDD VSS in[449] out[449] buffer
x_and449 VSS VDD in[449] clk out[449] AND2x2_ASAP7_75t_SRAM
x_buf450 VDD VSS in[450] out[450] buffer
x_and450 VSS VDD in[450] clk out[450] AND2x2_ASAP7_75t_SRAM
x_buf451 VDD VSS in[451] out[451] buffer
x_and451 VSS VDD in[451] clk out[451] AND2x2_ASAP7_75t_SRAM
x_buf452 VDD VSS in[452] out[452] buffer
x_and452 VSS VDD in[452] clk out[452] AND2x2_ASAP7_75t_SRAM
x_buf453 VDD VSS in[453] out[453] buffer
x_and453 VSS VDD in[453] clk out[453] AND2x2_ASAP7_75t_SRAM
x_buf454 VDD VSS in[454] out[454] buffer
x_and454 VSS VDD in[454] clk out[454] AND2x2_ASAP7_75t_SRAM
x_buf455 VDD VSS in[455] out[455] buffer
x_and455 VSS VDD in[455] clk out[455] AND2x2_ASAP7_75t_SRAM
x_buf456 VDD VSS in[456] out[456] buffer
x_and456 VSS VDD in[456] clk out[456] AND2x2_ASAP7_75t_SRAM
x_buf457 VDD VSS in[457] out[457] buffer
x_and457 VSS VDD in[457] clk out[457] AND2x2_ASAP7_75t_SRAM
x_buf458 VDD VSS in[458] out[458] buffer
x_and458 VSS VDD in[458] clk out[458] AND2x2_ASAP7_75t_SRAM
x_buf459 VDD VSS in[459] out[459] buffer
x_and459 VSS VDD in[459] clk out[459] AND2x2_ASAP7_75t_SRAM
x_buf460 VDD VSS in[460] out[460] buffer
x_and460 VSS VDD in[460] clk out[460] AND2x2_ASAP7_75t_SRAM
x_buf461 VDD VSS in[461] out[461] buffer
x_and461 VSS VDD in[461] clk out[461] AND2x2_ASAP7_75t_SRAM
x_buf462 VDD VSS in[462] out[462] buffer
x_and462 VSS VDD in[462] clk out[462] AND2x2_ASAP7_75t_SRAM
x_buf463 VDD VSS in[463] out[463] buffer
x_and463 VSS VDD in[463] clk out[463] AND2x2_ASAP7_75t_SRAM
x_buf464 VDD VSS in[464] out[464] buffer
x_and464 VSS VDD in[464] clk out[464] AND2x2_ASAP7_75t_SRAM
x_buf465 VDD VSS in[465] out[465] buffer
x_and465 VSS VDD in[465] clk out[465] AND2x2_ASAP7_75t_SRAM
x_buf466 VDD VSS in[466] out[466] buffer
x_and466 VSS VDD in[466] clk out[466] AND2x2_ASAP7_75t_SRAM
x_buf467 VDD VSS in[467] out[467] buffer
x_and467 VSS VDD in[467] clk out[467] AND2x2_ASAP7_75t_SRAM
x_buf468 VDD VSS in[468] out[468] buffer
x_and468 VSS VDD in[468] clk out[468] AND2x2_ASAP7_75t_SRAM
x_buf469 VDD VSS in[469] out[469] buffer
x_and469 VSS VDD in[469] clk out[469] AND2x2_ASAP7_75t_SRAM
x_buf470 VDD VSS in[470] out[470] buffer
x_and470 VSS VDD in[470] clk out[470] AND2x2_ASAP7_75t_SRAM
x_buf471 VDD VSS in[471] out[471] buffer
x_and471 VSS VDD in[471] clk out[471] AND2x2_ASAP7_75t_SRAM
x_buf472 VDD VSS in[472] out[472] buffer
x_and472 VSS VDD in[472] clk out[472] AND2x2_ASAP7_75t_SRAM
x_buf473 VDD VSS in[473] out[473] buffer
x_and473 VSS VDD in[473] clk out[473] AND2x2_ASAP7_75t_SRAM
x_buf474 VDD VSS in[474] out[474] buffer
x_and474 VSS VDD in[474] clk out[474] AND2x2_ASAP7_75t_SRAM
x_buf475 VDD VSS in[475] out[475] buffer
x_and475 VSS VDD in[475] clk out[475] AND2x2_ASAP7_75t_SRAM
x_buf476 VDD VSS in[476] out[476] buffer
x_and476 VSS VDD in[476] clk out[476] AND2x2_ASAP7_75t_SRAM
x_buf477 VDD VSS in[477] out[477] buffer
x_and477 VSS VDD in[477] clk out[477] AND2x2_ASAP7_75t_SRAM
x_buf478 VDD VSS in[478] out[478] buffer
x_and478 VSS VDD in[478] clk out[478] AND2x2_ASAP7_75t_SRAM
x_buf479 VDD VSS in[479] out[479] buffer
x_and479 VSS VDD in[479] clk out[479] AND2x2_ASAP7_75t_SRAM
x_buf480 VDD VSS in[480] out[480] buffer
x_and480 VSS VDD in[480] clk out[480] AND2x2_ASAP7_75t_SRAM
x_buf481 VDD VSS in[481] out[481] buffer
x_and481 VSS VDD in[481] clk out[481] AND2x2_ASAP7_75t_SRAM
x_buf482 VDD VSS in[482] out[482] buffer
x_and482 VSS VDD in[482] clk out[482] AND2x2_ASAP7_75t_SRAM
x_buf483 VDD VSS in[483] out[483] buffer
x_and483 VSS VDD in[483] clk out[483] AND2x2_ASAP7_75t_SRAM
x_buf484 VDD VSS in[484] out[484] buffer
x_and484 VSS VDD in[484] clk out[484] AND2x2_ASAP7_75t_SRAM
x_buf485 VDD VSS in[485] out[485] buffer
x_and485 VSS VDD in[485] clk out[485] AND2x2_ASAP7_75t_SRAM
x_buf486 VDD VSS in[486] out[486] buffer
x_and486 VSS VDD in[486] clk out[486] AND2x2_ASAP7_75t_SRAM
x_buf487 VDD VSS in[487] out[487] buffer
x_and487 VSS VDD in[487] clk out[487] AND2x2_ASAP7_75t_SRAM
x_buf488 VDD VSS in[488] out[488] buffer
x_and488 VSS VDD in[488] clk out[488] AND2x2_ASAP7_75t_SRAM
x_buf489 VDD VSS in[489] out[489] buffer
x_and489 VSS VDD in[489] clk out[489] AND2x2_ASAP7_75t_SRAM
x_buf490 VDD VSS in[490] out[490] buffer
x_and490 VSS VDD in[490] clk out[490] AND2x2_ASAP7_75t_SRAM
x_buf491 VDD VSS in[491] out[491] buffer
x_and491 VSS VDD in[491] clk out[491] AND2x2_ASAP7_75t_SRAM
x_buf492 VDD VSS in[492] out[492] buffer
x_and492 VSS VDD in[492] clk out[492] AND2x2_ASAP7_75t_SRAM
x_buf493 VDD VSS in[493] out[493] buffer
x_and493 VSS VDD in[493] clk out[493] AND2x2_ASAP7_75t_SRAM
x_buf494 VDD VSS in[494] out[494] buffer
x_and494 VSS VDD in[494] clk out[494] AND2x2_ASAP7_75t_SRAM
x_buf495 VDD VSS in[495] out[495] buffer
x_and495 VSS VDD in[495] clk out[495] AND2x2_ASAP7_75t_SRAM
x_buf496 VDD VSS in[496] out[496] buffer
x_and496 VSS VDD in[496] clk out[496] AND2x2_ASAP7_75t_SRAM
x_buf497 VDD VSS in[497] out[497] buffer
x_and497 VSS VDD in[497] clk out[497] AND2x2_ASAP7_75t_SRAM
x_buf498 VDD VSS in[498] out[498] buffer
x_and498 VSS VDD in[498] clk out[498] AND2x2_ASAP7_75t_SRAM
x_buf499 VDD VSS in[499] out[499] buffer
x_and499 VSS VDD in[499] clk out[499] AND2x2_ASAP7_75t_SRAM
x_buf500 VDD VSS in[500] out[500] buffer
x_and500 VSS VDD in[500] clk out[500] AND2x2_ASAP7_75t_SRAM
x_buf501 VDD VSS in[501] out[501] buffer
x_and501 VSS VDD in[501] clk out[501] AND2x2_ASAP7_75t_SRAM
x_buf502 VDD VSS in[502] out[502] buffer
x_and502 VSS VDD in[502] clk out[502] AND2x2_ASAP7_75t_SRAM
x_buf503 VDD VSS in[503] out[503] buffer
x_and503 VSS VDD in[503] clk out[503] AND2x2_ASAP7_75t_SRAM
x_buf504 VDD VSS in[504] out[504] buffer
x_and504 VSS VDD in[504] clk out[504] AND2x2_ASAP7_75t_SRAM
x_buf505 VDD VSS in[505] out[505] buffer
x_and505 VSS VDD in[505] clk out[505] AND2x2_ASAP7_75t_SRAM
x_buf506 VDD VSS in[506] out[506] buffer
x_and506 VSS VDD in[506] clk out[506] AND2x2_ASAP7_75t_SRAM
x_buf507 VDD VSS in[507] out[507] buffer
x_and507 VSS VDD in[507] clk out[507] AND2x2_ASAP7_75t_SRAM
x_buf508 VDD VSS in[508] out[508] buffer
x_and508 VSS VDD in[508] clk out[508] AND2x2_ASAP7_75t_SRAM
x_buf509 VDD VSS in[509] out[509] buffer
x_and509 VSS VDD in[509] clk out[509] AND2x2_ASAP7_75t_SRAM
x_buf510 VDD VSS in[510] out[510] buffer
x_and510 VSS VDD in[510] clk out[510] AND2x2_ASAP7_75t_SRAM
x_buf511 VDD VSS in[511] out[511] buffer
x_and511 VSS VDD in[511] clk out[511] AND2x2_ASAP7_75t_SRAM
.ends
.nodeset v(x_sram_arr0.x_cell0.q) = 0
.nodeset v(x_sram_arr0.x_cell1.q) = 0
.nodeset v(x_sram_arr0.x_cell2.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell3.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell4.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell5.q) = 0
.nodeset v(x_sram_arr0.x_cell6.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell7.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell8.q) = 0
.nodeset v(x_sram_arr0.x_cell9.q) = 0
.nodeset v(x_sram_arr0.x_cell10.q) = 0
.nodeset v(x_sram_arr0.x_cell11.q) = 0
.nodeset v(x_sram_arr0.x_cell12.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell13.q) = 0
.nodeset v(x_sram_arr0.x_cell14.q) = 0
.nodeset v(x_sram_arr0.x_cell15.q) = 0
.nodeset v(x_sram_arr0.x_cell16.q) = 0
.nodeset v(x_sram_arr0.x_cell17.q) = 0
.nodeset v(x_sram_arr0.x_cell18.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell19.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell20.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell21.q) = 0
.nodeset v(x_sram_arr0.x_cell22.q) = 0
.nodeset v(x_sram_arr0.x_cell23.q) = 0
.nodeset v(x_sram_arr0.x_cell24.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell25.q) = 0
.nodeset v(x_sram_arr0.x_cell26.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell27.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell28.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell29.q) = 0
.nodeset v(x_sram_arr0.x_cell30.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell31.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell32.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell33.q) = 0
.nodeset v(x_sram_arr0.x_cell34.q) = 0
.nodeset v(x_sram_arr0.x_cell35.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell36.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell37.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell38.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell39.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell40.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell41.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell42.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell43.q) = 0
.nodeset v(x_sram_arr0.x_cell44.q) = 0
.nodeset v(x_sram_arr0.x_cell45.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell46.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell47.q) = 0
.nodeset v(x_sram_arr0.x_cell48.q) = 0
.nodeset v(x_sram_arr0.x_cell49.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell50.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell51.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell52.q) = 0
.nodeset v(x_sram_arr0.x_cell53.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell54.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell55.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell56.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell57.q) = 0
.nodeset v(x_sram_arr0.x_cell58.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell59.q) = 0
.nodeset v(x_sram_arr0.x_cell60.q) = 0
.nodeset v(x_sram_arr0.x_cell61.q) = 0
.nodeset v(x_sram_arr0.x_cell62.q) = 0
.nodeset v(x_sram_arr0.x_cell63.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell64.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell65.q) = 0
.nodeset v(x_sram_arr0.x_cell66.q) = 0
.nodeset v(x_sram_arr0.x_cell67.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell68.q) = 0
.nodeset v(x_sram_arr0.x_cell69.q) = 0
.nodeset v(x_sram_arr0.x_cell70.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell71.q) = 0
.nodeset v(x_sram_arr0.x_cell72.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell73.q) = 0
.nodeset v(x_sram_arr0.x_cell74.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell75.q) = 0
.nodeset v(x_sram_arr0.x_cell76.q) = 0
.nodeset v(x_sram_arr0.x_cell77.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell78.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell79.q) = 0
.nodeset v(x_sram_arr0.x_cell80.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell81.q) = 0
.nodeset v(x_sram_arr0.x_cell82.q) = 0
.nodeset v(x_sram_arr0.x_cell83.q) = 0
.nodeset v(x_sram_arr0.x_cell84.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell85.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell86.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell87.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell88.q) = 0
.nodeset v(x_sram_arr0.x_cell89.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell90.q) = 0
.nodeset v(x_sram_arr0.x_cell91.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell92.q) = 0
.nodeset v(x_sram_arr0.x_cell93.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell94.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell95.q) = 0
.nodeset v(x_sram_arr0.x_cell96.q) = 0
.nodeset v(x_sram_arr0.x_cell97.q) = 0
.nodeset v(x_sram_arr0.x_cell98.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell99.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell100.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell101.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell102.q) = 0
.nodeset v(x_sram_arr0.x_cell103.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell104.q) = 0
.nodeset v(x_sram_arr0.x_cell105.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell106.q) = 0
.nodeset v(x_sram_arr0.x_cell107.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell108.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell109.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell110.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell111.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell112.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell113.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell114.q) = 0
.nodeset v(x_sram_arr0.x_cell115.q) = 0
.nodeset v(x_sram_arr0.x_cell116.q) = 0
.nodeset v(x_sram_arr0.x_cell117.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell118.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell119.q) = 0
.nodeset v(x_sram_arr0.x_cell120.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell121.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell122.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell123.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell124.q) = 0
.nodeset v(x_sram_arr0.x_cell125.q) = 0
.nodeset v(x_sram_arr0.x_cell126.q) = 0
.nodeset v(x_sram_arr0.x_cell127.q) = 0
.nodeset v(x_sram_arr0.x_cell128.q) = 0
.nodeset v(x_sram_arr0.x_cell129.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell130.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell131.q) = 0
.nodeset v(x_sram_arr0.x_cell132.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell133.q) = 0
.nodeset v(x_sram_arr0.x_cell134.q) = 0
.nodeset v(x_sram_arr0.x_cell135.q) = 0
.nodeset v(x_sram_arr0.x_cell136.q) = 0
.nodeset v(x_sram_arr0.x_cell137.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell138.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell139.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell140.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell141.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell142.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell143.q) = 0
.nodeset v(x_sram_arr0.x_cell144.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell145.q) = 0
.nodeset v(x_sram_arr0.x_cell146.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell147.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell148.q) = 0
.nodeset v(x_sram_arr0.x_cell149.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell150.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell151.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell152.q) = 0
.nodeset v(x_sram_arr0.x_cell153.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell154.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell155.q) = 0
.nodeset v(x_sram_arr0.x_cell156.q) = 0
.nodeset v(x_sram_arr0.x_cell157.q) = 0
.nodeset v(x_sram_arr0.x_cell158.q) = 0
.nodeset v(x_sram_arr0.x_cell159.q) = 0
.nodeset v(x_sram_arr0.x_cell160.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell161.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell162.q) = 0
.nodeset v(x_sram_arr0.x_cell163.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell164.q) = 0
.nodeset v(x_sram_arr0.x_cell165.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell166.q) = 0
.nodeset v(x_sram_arr0.x_cell167.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell168.q) = 0
.nodeset v(x_sram_arr0.x_cell169.q) = 0
.nodeset v(x_sram_arr0.x_cell170.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell171.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell172.q) = 0
.nodeset v(x_sram_arr0.x_cell173.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell174.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell175.q) = 0
.nodeset v(x_sram_arr0.x_cell176.q) = 0
.nodeset v(x_sram_arr0.x_cell177.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell178.q) = 0
.nodeset v(x_sram_arr0.x_cell179.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell180.q) = 0
.nodeset v(x_sram_arr0.x_cell181.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell182.q) = 0
.nodeset v(x_sram_arr0.x_cell183.q) = 0
.nodeset v(x_sram_arr0.x_cell184.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell185.q) = 0
.nodeset v(x_sram_arr0.x_cell186.q) = 0
.nodeset v(x_sram_arr0.x_cell187.q) = 0
.nodeset v(x_sram_arr0.x_cell188.q) = 0
.nodeset v(x_sram_arr0.x_cell189.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell190.q) = 0
.nodeset v(x_sram_arr0.x_cell191.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell192.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell193.q) = 0
.nodeset v(x_sram_arr0.x_cell194.q) = 0
.nodeset v(x_sram_arr0.x_cell195.q) = 0
.nodeset v(x_sram_arr0.x_cell196.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell197.q) = 0
.nodeset v(x_sram_arr0.x_cell198.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell199.q) = 0
.nodeset v(x_sram_arr0.x_cell200.q) = 0
.nodeset v(x_sram_arr0.x_cell201.q) = 0
.nodeset v(x_sram_arr0.x_cell202.q) = 0
.nodeset v(x_sram_arr0.x_cell203.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell204.q) = 0
.nodeset v(x_sram_arr0.x_cell205.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell206.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell207.q) = 0
.nodeset v(x_sram_arr0.x_cell208.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell209.q) = 0
.nodeset v(x_sram_arr0.x_cell210.q) = 0
.nodeset v(x_sram_arr0.x_cell211.q) = 0
.nodeset v(x_sram_arr0.x_cell212.q) = 0
.nodeset v(x_sram_arr0.x_cell213.q) = 0
.nodeset v(x_sram_arr0.x_cell214.q) = 0
.nodeset v(x_sram_arr0.x_cell215.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell216.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell217.q) = 0
.nodeset v(x_sram_arr0.x_cell218.q) = 0
.nodeset v(x_sram_arr0.x_cell219.q) = 0
.nodeset v(x_sram_arr0.x_cell220.q) = 0
.nodeset v(x_sram_arr0.x_cell221.q) = 0
.nodeset v(x_sram_arr0.x_cell222.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell223.q) = 0
.nodeset v(x_sram_arr0.x_cell224.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell225.q) = 0
.nodeset v(x_sram_arr0.x_cell226.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell227.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell228.q) = 0
.nodeset v(x_sram_arr0.x_cell229.q) = 0
.nodeset v(x_sram_arr0.x_cell230.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell231.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell232.q) = 0
.nodeset v(x_sram_arr0.x_cell233.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell234.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell235.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell236.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell237.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell238.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell239.q) = 0
.nodeset v(x_sram_arr0.x_cell240.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell241.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell242.q) = 0
.nodeset v(x_sram_arr0.x_cell243.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell244.q) = 0
.nodeset v(x_sram_arr0.x_cell245.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell246.q) = 0
.nodeset v(x_sram_arr0.x_cell247.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell248.q) = 0
.nodeset v(x_sram_arr0.x_cell249.q) = 0
.nodeset v(x_sram_arr0.x_cell250.q) = 0
.nodeset v(x_sram_arr0.x_cell251.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell252.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell253.q) = 0
.nodeset v(x_sram_arr0.x_cell254.q) = 0
.nodeset v(x_sram_arr0.x_cell255.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell256.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell257.q) = 0
.nodeset v(x_sram_arr0.x_cell258.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell259.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell260.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell261.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell262.q) = 0
.nodeset v(x_sram_arr0.x_cell263.q) = 0
.nodeset v(x_sram_arr0.x_cell264.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell265.q) = 0
.nodeset v(x_sram_arr0.x_cell266.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell267.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell268.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell269.q) = 0
.nodeset v(x_sram_arr0.x_cell270.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell271.q) = 0
.nodeset v(x_sram_arr0.x_cell272.q) = 0
.nodeset v(x_sram_arr0.x_cell273.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell274.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell275.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell276.q) = 0
.nodeset v(x_sram_arr0.x_cell277.q) = 0
.nodeset v(x_sram_arr0.x_cell278.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell279.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell280.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell281.q) = 0
.nodeset v(x_sram_arr0.x_cell282.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell283.q) = 0
.nodeset v(x_sram_arr0.x_cell284.q) = 0
.nodeset v(x_sram_arr0.x_cell285.q) = 0
.nodeset v(x_sram_arr0.x_cell286.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell287.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell288.q) = 0
.nodeset v(x_sram_arr0.x_cell289.q) = 0
.nodeset v(x_sram_arr0.x_cell290.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell291.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell292.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell293.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell294.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell295.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell296.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell297.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell298.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell299.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell300.q) = 0
.nodeset v(x_sram_arr0.x_cell301.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell302.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell303.q) = 0
.nodeset v(x_sram_arr0.x_cell304.q) = 0
.nodeset v(x_sram_arr0.x_cell305.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell306.q) = 0
.nodeset v(x_sram_arr0.x_cell307.q) = 0
.nodeset v(x_sram_arr0.x_cell308.q) = 0
.nodeset v(x_sram_arr0.x_cell309.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell310.q) = 0
.nodeset v(x_sram_arr0.x_cell311.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell312.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell313.q) = 0
.nodeset v(x_sram_arr0.x_cell314.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell315.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell316.q) = 0
.nodeset v(x_sram_arr0.x_cell317.q) = 0
.nodeset v(x_sram_arr0.x_cell318.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell319.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell320.q) = 0
.nodeset v(x_sram_arr0.x_cell321.q) = 0
.nodeset v(x_sram_arr0.x_cell322.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell323.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell324.q) = 0
.nodeset v(x_sram_arr0.x_cell325.q) = 0
.nodeset v(x_sram_arr0.x_cell326.q) = 0
.nodeset v(x_sram_arr0.x_cell327.q) = 0
.nodeset v(x_sram_arr0.x_cell328.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell329.q) = 0
.nodeset v(x_sram_arr0.x_cell330.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell331.q) = 0
.nodeset v(x_sram_arr0.x_cell332.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell333.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell334.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell335.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell336.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell337.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell338.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell339.q) = 0
.nodeset v(x_sram_arr0.x_cell340.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell341.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell342.q) = 0
.nodeset v(x_sram_arr0.x_cell343.q) = 0
.nodeset v(x_sram_arr0.x_cell344.q) = 0
.nodeset v(x_sram_arr0.x_cell345.q) = 0
.nodeset v(x_sram_arr0.x_cell346.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell347.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell348.q) = 0
.nodeset v(x_sram_arr0.x_cell349.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell350.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell351.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell352.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell353.q) = 0
.nodeset v(x_sram_arr0.x_cell354.q) = 0
.nodeset v(x_sram_arr0.x_cell355.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell356.q) = 0
.nodeset v(x_sram_arr0.x_cell357.q) = 0
.nodeset v(x_sram_arr0.x_cell358.q) = 0
.nodeset v(x_sram_arr0.x_cell359.q) = 0
.nodeset v(x_sram_arr0.x_cell360.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell361.q) = 0
.nodeset v(x_sram_arr0.x_cell362.q) = 0
.nodeset v(x_sram_arr0.x_cell363.q) = 0
.nodeset v(x_sram_arr0.x_cell364.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell365.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell366.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell367.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell368.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell369.q) = 0
.nodeset v(x_sram_arr0.x_cell370.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell371.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell372.q) = 0
.nodeset v(x_sram_arr0.x_cell373.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell374.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell375.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell376.q) = 0
.nodeset v(x_sram_arr0.x_cell377.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell378.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell379.q) = 0
.nodeset v(x_sram_arr0.x_cell380.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell381.q) = 0
.nodeset v(x_sram_arr0.x_cell382.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell383.q) = 0
.nodeset v(x_sram_arr0.x_cell384.q) = 0
.nodeset v(x_sram_arr0.x_cell385.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell386.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell387.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell388.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell389.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell390.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell391.q) = 0
.nodeset v(x_sram_arr0.x_cell392.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell393.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell394.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell395.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell396.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell397.q) = 0
.nodeset v(x_sram_arr0.x_cell398.q) = 0
.nodeset v(x_sram_arr0.x_cell399.q) = 0
.nodeset v(x_sram_arr0.x_cell400.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell401.q) = 0
.nodeset v(x_sram_arr0.x_cell402.q) = 0
.nodeset v(x_sram_arr0.x_cell403.q) = 0
.nodeset v(x_sram_arr0.x_cell404.q) = 0
.nodeset v(x_sram_arr0.x_cell405.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell406.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell407.q) = 0
.nodeset v(x_sram_arr0.x_cell408.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell409.q) = 0
.nodeset v(x_sram_arr0.x_cell410.q) = 0
.nodeset v(x_sram_arr0.x_cell411.q) = 0
.nodeset v(x_sram_arr0.x_cell412.q) = 0
.nodeset v(x_sram_arr0.x_cell413.q) = 0
.nodeset v(x_sram_arr0.x_cell414.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell415.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell416.q) = 0
.nodeset v(x_sram_arr0.x_cell417.q) = 0
.nodeset v(x_sram_arr0.x_cell418.q) = 0
.nodeset v(x_sram_arr0.x_cell419.q) = 0
.nodeset v(x_sram_arr0.x_cell420.q) = 0
.nodeset v(x_sram_arr0.x_cell421.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell422.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell423.q) = 0
.nodeset v(x_sram_arr0.x_cell424.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell425.q) = 0
.nodeset v(x_sram_arr0.x_cell426.q) = 0
.nodeset v(x_sram_arr0.x_cell427.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell428.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell429.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell430.q) = 0
.nodeset v(x_sram_arr0.x_cell431.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell432.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell433.q) = 0
.nodeset v(x_sram_arr0.x_cell434.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell435.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell436.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell437.q) = 0
.nodeset v(x_sram_arr0.x_cell438.q) = 0
.nodeset v(x_sram_arr0.x_cell439.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell440.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell441.q) = 0
.nodeset v(x_sram_arr0.x_cell442.q) = 0
.nodeset v(x_sram_arr0.x_cell443.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell444.q) = 0
.nodeset v(x_sram_arr0.x_cell445.q) = 0
.nodeset v(x_sram_arr0.x_cell446.q) = 0
.nodeset v(x_sram_arr0.x_cell447.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell448.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell449.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell450.q) = 0
.nodeset v(x_sram_arr0.x_cell451.q) = 0
.nodeset v(x_sram_arr0.x_cell452.q) = 0
.nodeset v(x_sram_arr0.x_cell453.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell454.q) = 0
.nodeset v(x_sram_arr0.x_cell455.q) = 0
.nodeset v(x_sram_arr0.x_cell456.q) = 0
.nodeset v(x_sram_arr0.x_cell457.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell458.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell459.q) = 0
.nodeset v(x_sram_arr0.x_cell460.q) = 0
.nodeset v(x_sram_arr0.x_cell461.q) = 0
.nodeset v(x_sram_arr0.x_cell462.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell463.q) = 0
.nodeset v(x_sram_arr0.x_cell464.q) = 0
.nodeset v(x_sram_arr0.x_cell465.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell466.q) = 0
.nodeset v(x_sram_arr0.x_cell467.q) = 0
.nodeset v(x_sram_arr0.x_cell468.q) = 0
.nodeset v(x_sram_arr0.x_cell469.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell470.q) = 0
.nodeset v(x_sram_arr0.x_cell471.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell472.q) = 0
.nodeset v(x_sram_arr0.x_cell473.q) = 0
.nodeset v(x_sram_arr0.x_cell474.q) = 0
.nodeset v(x_sram_arr0.x_cell475.q) = 0
.nodeset v(x_sram_arr0.x_cell476.q) = 0
.nodeset v(x_sram_arr0.x_cell477.q) = 0
.nodeset v(x_sram_arr0.x_cell478.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell479.q) = 0
.nodeset v(x_sram_arr0.x_cell480.q) = 0
.nodeset v(x_sram_arr0.x_cell481.q) = 0
.nodeset v(x_sram_arr0.x_cell482.q) = 0
.nodeset v(x_sram_arr0.x_cell483.q) = 0
.nodeset v(x_sram_arr0.x_cell484.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell485.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell486.q) = 0
.nodeset v(x_sram_arr0.x_cell487.q) = 0
.nodeset v(x_sram_arr0.x_cell488.q) = 0
.nodeset v(x_sram_arr0.x_cell489.q) = 0
.nodeset v(x_sram_arr0.x_cell490.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell491.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell492.q) = 0
.nodeset v(x_sram_arr0.x_cell493.q) = 0
.nodeset v(x_sram_arr0.x_cell494.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell495.q) = 0
.nodeset v(x_sram_arr0.x_cell496.q) = 0
.nodeset v(x_sram_arr0.x_cell497.q) = 0
.nodeset v(x_sram_arr0.x_cell498.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell499.q) = 0
.nodeset v(x_sram_arr0.x_cell500.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell501.q) = 0
.nodeset v(x_sram_arr0.x_cell502.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell503.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell504.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell505.q) = 0
.nodeset v(x_sram_arr0.x_cell506.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell507.q) = 0
.nodeset v(x_sram_arr0.x_cell508.q) = v_vdd
.nodeset v(x_sram_arr0.x_cell509.q) = 0
.nodeset v(x_sram_arr0.x_cell510.q) = 0
.nodeset v(x_sram_arr0.x_cell511.q) = 0
