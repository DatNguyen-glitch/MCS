.SUBCKT decoder_6to64 VDD VSS  clk rst_n in_addr[5] in_addr[4] in_addr[3] in_addr[2] in_addr[1] in_addr[0] wordline[63] wordline[62] wordline[61] wordline[60] wordline[59] wordline[58] wordline[57] wordline[56] wordline[55] wordline[54] wordline[53] wordline[52] wordline[51] wordline[50] wordline[49] wordline[48] wordline[47] wordline[46] wordline[45] wordline[44] wordline[43] wordline[42] wordline[41] wordline[40] wordline[39] wordline[38] wordline[37] wordline[36] wordline[35] wordline[34] wordline[33] wordline[32] wordline[31] wordline[30] wordline[29] wordline[28] wordline[27] wordline[26] wordline[25] wordline[24] wordline[23] wordline[22] wordline[21] wordline[20] wordline[19] wordline[18] wordline[17] wordline[16] wordline[15] wordline[14] wordline[13] wordline[12] wordline[11] wordline[10] wordline[9] wordline[8] wordline[7] wordline[6] wordline[5] wordline[4] wordline[3] wordline[2] wordline[1] wordline[0]
Xmsb_decoder addr[5] addr[4] addr[3] msb_en[7] msb_en[6] msb_en[5] msb_en[4] msb_en[3] msb_en[2] msb_en[1] VDD VSS  msb_en[0] decoder_3to8_8
Xlsb_decoder_group_0__lsb_decoder n17 n16 n15 lsb_decoder_group_0__lsb_out[7] lsb_decoder_group_0__lsb_out[6] lsb_decoder_group_0__lsb_out[5] lsb_decoder_group_0__lsb_out[4] lsb_decoder_group_0__lsb_out[3] lsb_decoder_group_0__lsb_out[2] lsb_decoder_group_0__lsb_out[1] VDD VSS  lsb_decoder_group_0__lsb_out[0] decoder_3to8_7
Xlsb_decoder_group_1__lsb_decoder n17 n16 n15 lsb_decoder_group_1__lsb_out[7] lsb_decoder_group_1__lsb_out[6] lsb_decoder_group_1__lsb_out[5] lsb_decoder_group_1__lsb_out[4] lsb_decoder_group_1__lsb_out[3] lsb_decoder_group_1__lsb_out[2] lsb_decoder_group_1__lsb_out[1] VDD VSS  lsb_decoder_group_1__lsb_out[0] decoder_3to8_6
Xlsb_decoder_group_2__lsb_decoder n17 n16 n15 lsb_decoder_group_2__lsb_out[7] lsb_decoder_group_2__lsb_out[6] lsb_decoder_group_2__lsb_out[5] lsb_decoder_group_2__lsb_out[4] lsb_decoder_group_2__lsb_out[3] lsb_decoder_group_2__lsb_out[2] lsb_decoder_group_2__lsb_out[1] VDD VSS  lsb_decoder_group_2__lsb_out[0] decoder_3to8_5
Xlsb_decoder_group_3__lsb_decoder n17 n16 n15 lsb_decoder_group_3__lsb_out[7] lsb_decoder_group_3__lsb_out[6] lsb_decoder_group_3__lsb_out[5] lsb_decoder_group_3__lsb_out[4] lsb_decoder_group_3__lsb_out[3] lsb_decoder_group_3__lsb_out[2] lsb_decoder_group_3__lsb_out[1] VDD VSS  lsb_decoder_group_3__lsb_out[0] decoder_3to8_4
Xlsb_decoder_group_4__lsb_decoder n17 n16 n15 lsb_decoder_group_4__lsb_out[7] lsb_decoder_group_4__lsb_out[6] lsb_decoder_group_4__lsb_out[5] lsb_decoder_group_4__lsb_out[4] lsb_decoder_group_4__lsb_out[3] lsb_decoder_group_4__lsb_out[2] lsb_decoder_group_4__lsb_out[1] VDD VSS  lsb_decoder_group_4__lsb_out[0] decoder_3to8_3
Xlsb_decoder_group_5__lsb_decoder n17 n16 n15 lsb_decoder_group_5__lsb_out[7] lsb_decoder_group_5__lsb_out[6] lsb_decoder_group_5__lsb_out[5] lsb_decoder_group_5__lsb_out[4] lsb_decoder_group_5__lsb_out[3] lsb_decoder_group_5__lsb_out[2] lsb_decoder_group_5__lsb_out[1] VDD VSS  lsb_decoder_group_5__lsb_out[0] decoder_3to8_2
Xlsb_decoder_group_6__lsb_decoder n17 n16 n15 lsb_decoder_group_6__lsb_out[7] lsb_decoder_group_6__lsb_out[6] lsb_decoder_group_6__lsb_out[5] lsb_decoder_group_6__lsb_out[4] lsb_decoder_group_6__lsb_out[3] lsb_decoder_group_6__lsb_out[2] lsb_decoder_group_6__lsb_out[1] VDD VSS  lsb_decoder_group_6__lsb_out[0] decoder_3to8_1
Xlsb_decoder_group_7__lsb_decoder n17 n16 n15 lsb_decoder_group_7__lsb_out[7] lsb_decoder_group_7__lsb_out[6] lsb_decoder_group_7__lsb_out[5] lsb_decoder_group_7__lsb_out[4] lsb_decoder_group_7__lsb_out[3] lsb_decoder_group_7__lsb_out[2] lsb_decoder_group_7__lsb_out[1] VDD VSS  lsb_decoder_group_7__lsb_out[0] decoder_3to8_0
XU3 in_addr[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU5 in_addr[1] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
XU7 in_addr[2] VDD VSS  n5 INVx1_ASAP7_75t_SRAM
XU9 in_addr[3] VDD VSS  n7 INVx1_ASAP7_75t_SRAM
XU11 in_addr[4] VDD VSS  n9 INVx1_ASAP7_75t_SRAM
XU13 in_addr[5] VDD VSS  n11 INVx1_ASAP7_75t_SRAM
XU15 rst_n VDD VSS  n13 INVx1_ASAP7_75t_SRAM
XU16 lsb_decoder_group_1__lsb_out[1] msb_en[1] VDD VSS  wordline[9] OR2x2_ASAP7_75t_SRAM
XU17 lsb_decoder_group_1__lsb_out[0] msb_en[1] VDD VSS  wordline[8] OR2x2_ASAP7_75t_SRAM
XU18 lsb_decoder_group_0__lsb_out[7] msb_en[0] VDD VSS  wordline[7] OR2x2_ASAP7_75t_SRAM
XU19 lsb_decoder_group_0__lsb_out[6] msb_en[0] VDD VSS  wordline[6] OR2x2_ASAP7_75t_SRAM
XU20 lsb_decoder_group_7__lsb_out[7] msb_en[7] VDD VSS  wordline[63] OR2x2_ASAP7_75t_SRAM
XU21 lsb_decoder_group_7__lsb_out[6] msb_en[7] VDD VSS  wordline[62] OR2x2_ASAP7_75t_SRAM
XU22 lsb_decoder_group_7__lsb_out[5] msb_en[7] VDD VSS  wordline[61] OR2x2_ASAP7_75t_SRAM
XU23 lsb_decoder_group_7__lsb_out[4] msb_en[7] VDD VSS  wordline[60] OR2x2_ASAP7_75t_SRAM
XU24 lsb_decoder_group_0__lsb_out[5] msb_en[0] VDD VSS  wordline[5] OR2x2_ASAP7_75t_SRAM
XU25 lsb_decoder_group_7__lsb_out[3] msb_en[7] VDD VSS  wordline[59] OR2x2_ASAP7_75t_SRAM
XU26 lsb_decoder_group_7__lsb_out[2] msb_en[7] VDD VSS  wordline[58] OR2x2_ASAP7_75t_SRAM
XU27 lsb_decoder_group_7__lsb_out[1] msb_en[7] VDD VSS  wordline[57] OR2x2_ASAP7_75t_SRAM
XU28 lsb_decoder_group_7__lsb_out[0] msb_en[7] VDD VSS  wordline[56] OR2x2_ASAP7_75t_SRAM
XU29 lsb_decoder_group_6__lsb_out[7] msb_en[6] VDD VSS  wordline[55] OR2x2_ASAP7_75t_SRAM
XU30 lsb_decoder_group_6__lsb_out[6] msb_en[6] VDD VSS  wordline[54] OR2x2_ASAP7_75t_SRAM
XU31 lsb_decoder_group_6__lsb_out[5] msb_en[6] VDD VSS  wordline[53] OR2x2_ASAP7_75t_SRAM
XU32 lsb_decoder_group_6__lsb_out[4] msb_en[6] VDD VSS  wordline[52] OR2x2_ASAP7_75t_SRAM
XU33 lsb_decoder_group_6__lsb_out[3] msb_en[6] VDD VSS  wordline[51] OR2x2_ASAP7_75t_SRAM
XU34 lsb_decoder_group_6__lsb_out[2] msb_en[6] VDD VSS  wordline[50] OR2x2_ASAP7_75t_SRAM
XU35 lsb_decoder_group_0__lsb_out[4] msb_en[0] VDD VSS  wordline[4] OR2x2_ASAP7_75t_SRAM
XU36 lsb_decoder_group_6__lsb_out[1] msb_en[6] VDD VSS  wordline[49] OR2x2_ASAP7_75t_SRAM
XU37 lsb_decoder_group_6__lsb_out[0] msb_en[6] VDD VSS  wordline[48] OR2x2_ASAP7_75t_SRAM
XU38 lsb_decoder_group_5__lsb_out[7] msb_en[5] VDD VSS  wordline[47] OR2x2_ASAP7_75t_SRAM
XU39 lsb_decoder_group_5__lsb_out[6] msb_en[5] VDD VSS  wordline[46] OR2x2_ASAP7_75t_SRAM
XU40 lsb_decoder_group_5__lsb_out[5] msb_en[5] VDD VSS  wordline[45] OR2x2_ASAP7_75t_SRAM
XU41 lsb_decoder_group_5__lsb_out[4] msb_en[5] VDD VSS  wordline[44] OR2x2_ASAP7_75t_SRAM
XU42 lsb_decoder_group_5__lsb_out[3] msb_en[5] VDD VSS  wordline[43] OR2x2_ASAP7_75t_SRAM
XU43 lsb_decoder_group_5__lsb_out[2] msb_en[5] VDD VSS  wordline[42] OR2x2_ASAP7_75t_SRAM
XU44 lsb_decoder_group_5__lsb_out[1] msb_en[5] VDD VSS  wordline[41] OR2x2_ASAP7_75t_SRAM
XU45 lsb_decoder_group_5__lsb_out[0] msb_en[5] VDD VSS  wordline[40] OR2x2_ASAP7_75t_SRAM
XU46 lsb_decoder_group_0__lsb_out[3] msb_en[0] VDD VSS  wordline[3] OR2x2_ASAP7_75t_SRAM
XU47 lsb_decoder_group_4__lsb_out[7] msb_en[4] VDD VSS  wordline[39] OR2x2_ASAP7_75t_SRAM
XU48 lsb_decoder_group_4__lsb_out[6] msb_en[4] VDD VSS  wordline[38] OR2x2_ASAP7_75t_SRAM
XU49 lsb_decoder_group_4__lsb_out[5] msb_en[4] VDD VSS  wordline[37] OR2x2_ASAP7_75t_SRAM
XU50 lsb_decoder_group_4__lsb_out[4] msb_en[4] VDD VSS  wordline[36] OR2x2_ASAP7_75t_SRAM
XU51 lsb_decoder_group_4__lsb_out[3] msb_en[4] VDD VSS  wordline[35] OR2x2_ASAP7_75t_SRAM
XU52 lsb_decoder_group_4__lsb_out[2] msb_en[4] VDD VSS  wordline[34] OR2x2_ASAP7_75t_SRAM
XU53 lsb_decoder_group_4__lsb_out[1] msb_en[4] VDD VSS  wordline[33] OR2x2_ASAP7_75t_SRAM
XU54 lsb_decoder_group_4__lsb_out[0] msb_en[4] VDD VSS  wordline[32] OR2x2_ASAP7_75t_SRAM
XU55 lsb_decoder_group_3__lsb_out[7] msb_en[3] VDD VSS  wordline[31] OR2x2_ASAP7_75t_SRAM
XU56 lsb_decoder_group_3__lsb_out[6] msb_en[3] VDD VSS  wordline[30] OR2x2_ASAP7_75t_SRAM
XU57 lsb_decoder_group_0__lsb_out[2] msb_en[0] VDD VSS  wordline[2] OR2x2_ASAP7_75t_SRAM
XU58 lsb_decoder_group_3__lsb_out[5] msb_en[3] VDD VSS  wordline[29] OR2x2_ASAP7_75t_SRAM
XU59 lsb_decoder_group_3__lsb_out[4] msb_en[3] VDD VSS  wordline[28] OR2x2_ASAP7_75t_SRAM
XU60 lsb_decoder_group_3__lsb_out[3] msb_en[3] VDD VSS  wordline[27] OR2x2_ASAP7_75t_SRAM
XU61 lsb_decoder_group_3__lsb_out[2] msb_en[3] VDD VSS  wordline[26] OR2x2_ASAP7_75t_SRAM
XU62 lsb_decoder_group_3__lsb_out[1] msb_en[3] VDD VSS  wordline[25] OR2x2_ASAP7_75t_SRAM
XU63 lsb_decoder_group_3__lsb_out[0] msb_en[3] VDD VSS  wordline[24] OR2x2_ASAP7_75t_SRAM
XU64 lsb_decoder_group_2__lsb_out[7] msb_en[2] VDD VSS  wordline[23] OR2x2_ASAP7_75t_SRAM
XU65 lsb_decoder_group_2__lsb_out[6] msb_en[2] VDD VSS  wordline[22] OR2x2_ASAP7_75t_SRAM
XU66 lsb_decoder_group_2__lsb_out[5] msb_en[2] VDD VSS  wordline[21] OR2x2_ASAP7_75t_SRAM
XU67 lsb_decoder_group_2__lsb_out[4] msb_en[2] VDD VSS  wordline[20] OR2x2_ASAP7_75t_SRAM
XU68 lsb_decoder_group_0__lsb_out[1] msb_en[0] VDD VSS  wordline[1] OR2x2_ASAP7_75t_SRAM
XU69 lsb_decoder_group_2__lsb_out[3] msb_en[2] VDD VSS  wordline[19] OR2x2_ASAP7_75t_SRAM
XU70 lsb_decoder_group_2__lsb_out[2] msb_en[2] VDD VSS  wordline[18] OR2x2_ASAP7_75t_SRAM
XU71 lsb_decoder_group_2__lsb_out[1] msb_en[2] VDD VSS  wordline[17] OR2x2_ASAP7_75t_SRAM
XU72 lsb_decoder_group_2__lsb_out[0] msb_en[2] VDD VSS  wordline[16] OR2x2_ASAP7_75t_SRAM
XU73 lsb_decoder_group_1__lsb_out[7] msb_en[1] VDD VSS  wordline[15] OR2x2_ASAP7_75t_SRAM
XU74 lsb_decoder_group_1__lsb_out[6] msb_en[1] VDD VSS  wordline[14] OR2x2_ASAP7_75t_SRAM
XU75 lsb_decoder_group_1__lsb_out[5] msb_en[1] VDD VSS  wordline[13] OR2x2_ASAP7_75t_SRAM
XU76 lsb_decoder_group_1__lsb_out[4] msb_en[1] VDD VSS  wordline[12] OR2x2_ASAP7_75t_SRAM
XU77 lsb_decoder_group_1__lsb_out[3] msb_en[1] VDD VSS  wordline[11] OR2x2_ASAP7_75t_SRAM
XU78 lsb_decoder_group_1__lsb_out[2] msb_en[1] VDD VSS  wordline[10] OR2x2_ASAP7_75t_SRAM
XU79 lsb_decoder_group_0__lsb_out[0] msb_en[0] VDD VSS  wordline[0] OR2x2_ASAP7_75t_SRAM
Xaddr_reg_5_ n11 clk n13 n14 VDD VSS  addr[5] ASYNC_DFFHx1_ASAP7_75t_SRAM
Xaddr_reg_4_ n9 clk n13 n14 VDD VSS  addr[4] ASYNC_DFFHx1_ASAP7_75t_SRAM
Xaddr_reg_3_ n7 clk n13 n14 VDD VSS  addr[3] ASYNC_DFFHx1_ASAP7_75t_SRAM
Xaddr_reg_2_ n5 clk n13 n14 VDD VSS  addr[2] ASYNC_DFFHx1_ASAP7_75t_SRAM
Xaddr_reg_1_ n3 clk n13 n14 VDD VSS  addr[1] ASYNC_DFFHx1_ASAP7_75t_SRAM
Xaddr_reg_0_ n1 clk n13 n14 VDD VSS  addr[0] ASYNC_DFFHx1_ASAP7_75t_SRAM
XU80 VDD VSS  n14 TIELOx1_ASAP7_75t_SRAM
XU81 addr[0] VDD VSS  n15 HB1xp67_ASAP7_75t_SRAM
XU82 addr[1] VDD VSS  n16 HB1xp67_ASAP7_75t_SRAM
XU83 addr[2] VDD VSS  n17 HB1xp67_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_7 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_6 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_5 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_4 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_3 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_2 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_1 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_0 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n1 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n1 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n3 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n1 n3 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n3 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n3 n1 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
XU1 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU2 a[0] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU3 a[2] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
.ENDS


.SUBCKT decoder_3to8_8 a[2] a[1] a[0] word[7] word[6] word[5] word[4] word[3] word[2] VDD VSS  word[1] word[0]
XU1 a[2] VDD VSS  n1 INVx1_ASAP7_75t_SRAM
XU2 a[1] VDD VSS  n2 INVx1_ASAP7_75t_SRAM
XU3 a[0] VDD VSS  n3 INVx1_ASAP7_75t_SRAM
XU4 a[1] a[0] a[2] VDD VSS  word[7] NAND3xp33_ASAP7_75t_SRAM
XU5 a[1] n3 a[2] VDD VSS  word[6] NAND3xp33_ASAP7_75t_SRAM
XU6 a[0] n2 a[2] VDD VSS  word[5] NAND3xp33_ASAP7_75t_SRAM
XU7 n3 n2 a[2] VDD VSS  word[4] NAND3xp33_ASAP7_75t_SRAM
XU8 a[0] n1 a[1] VDD VSS  word[3] NAND3xp33_ASAP7_75t_SRAM
XU9 n3 n1 a[1] VDD VSS  word[2] NAND3xp33_ASAP7_75t_SRAM
XU10 n2 n1 a[0] VDD VSS  word[1] NAND3xp33_ASAP7_75t_SRAM
XU11 n2 n1 n3 VDD VSS  word[0] NAND3xp33_ASAP7_75t_SRAM
.ENDS


