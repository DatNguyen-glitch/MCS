.SUBCKT decoder_6to64 clk in_addr[5] in_addr[4] in_addr[3] in_addr[2] in_addr[1] in_addr[0] wordline[63] wordline[62] wordline[61] wordline[60] wordline[59] wordline[58] wordline[57] wordline[56] wordline[55] wordline[54] wordline[53] wordline[52] wordline[51] wordline[50] wordline[49] wordline[48] wordline[47] wordline[46] wordline[45] wordline[44] wordline[43] wordline[42] wordline[41] wordline[40] wordline[39] wordline[38] wordline[37] wordline[36] wordline[35] wordline[34] wordline[33] wordline[32] wordline[31] wordline[30] wordline[29] wordline[28] wordline[27] wordline[26] wordline[25] wordline[24] wordline[23] wordline[22] wordline[21] wordline[20] wordline[19] wordline[18] wordline[17] wordline[16] wordline[15] wordline[14] wordline[13] wordline[12] wordline[11] wordline[10] wordline[9] wordline[8] wordline[7] wordline[6] wordline[5] wordline[4] wordline[3] wordline[2] wordline[1] wordline[0]
XU90 clk n46 INVx4_ASAP7_75t_SRAM
XU91 in_addr[0] n24 INVx5_ASAP7_75t_SRAM
XU92 in_addr[3] n25 INVx5_ASAP7_75t_SRAM
XU93 in_addr[4] n26 INVx5_ASAP7_75t_SRAM
XU94 in_addr[5] n27 INVx5_ASAP7_75t_SRAM
XU95 in_addr[1] n28 INVx5_ASAP7_75t_SRAM
XU96 in_addr[3] n29 INVx5_ASAP7_75t_SRAM
XU97 in_addr[3] n30 INVx5_ASAP7_75t_SRAM
XU98 in_addr[3] n39 INVx5_ASAP7_75t_SRAM
XU99 in_addr[0] n31 INVx5_ASAP7_75t_SRAM
XU100 in_addr[0] n32 INVx5_ASAP7_75t_SRAM
XU101 in_addr[4] n33 INVx5_ASAP7_75t_SRAM
XU102 in_addr[4] n34 INVx5_ASAP7_75t_SRAM
XU103 in_addr[0] n49 INVx5_ASAP7_75t_SRAM
XU104 in_addr[4] n40 INVx5_ASAP7_75t_SRAM
XU105 n61 n43 wordline[6] NOR2xp67_ASAP7_75t_SRAM
XU106 n61 n45 wordline[5] NOR2xp67_ASAP7_75t_SRAM
XU107 n61 n44 wordline[4] NOR2xp67_ASAP7_75t_SRAM
XU108 n42 n51 wordline[55] NOR2xp67_ASAP7_75t_SRAM
XU109 n42 n55 wordline[47] NOR2xp67_ASAP7_75t_SRAM
XU110 n42 n56 wordline[39] NOR2xp67_ASAP7_75t_SRAM
XU111 n42 n52 wordline[23] NOR2xp67_ASAP7_75t_SRAM
XU112 n42 n53 wordline[15] NOR2xp67_ASAP7_75t_SRAM
XU113 n42 n57 wordline[31] NOR2xp67_ASAP7_75t_SRAM
XU114 n61 n42 wordline[7] NOR2xp67_ASAP7_75t_SRAM
XU115 n43 n57 wordline[30] NOR2xp67_ASAP7_75t_SRAM
XU116 n43 n53 wordline[14] NOR2xp67_ASAP7_75t_SRAM
XU117 n43 n55 wordline[46] NOR2xp67_ASAP7_75t_SRAM
XU118 n43 n52 wordline[22] NOR2xp67_ASAP7_75t_SRAM
XU119 n43 n54 wordline[62] NOR2xp67_ASAP7_75t_SRAM
XU120 n43 n56 wordline[38] NOR2xp67_ASAP7_75t_SRAM
XU121 n44 n53 wordline[12] NOR2xp67_ASAP7_75t_SRAM
XU122 n44 n52 wordline[20] NOR2xp67_ASAP7_75t_SRAM
XU123 n44 n57 wordline[28] NOR2xp67_ASAP7_75t_SRAM
XU124 n44 n51 wordline[52] NOR2xp67_ASAP7_75t_SRAM
XU125 n44 n55 wordline[44] NOR2xp67_ASAP7_75t_SRAM
XU126 n45 n51 wordline[53] NOR2xp67_ASAP7_75t_SRAM
XU127 n44 n54 wordline[60] NOR2xp67_ASAP7_75t_SRAM
XU128 n44 n56 wordline[36] NOR2xp67_ASAP7_75t_SRAM
XU129 n45 n55 wordline[45] NOR2xp67_ASAP7_75t_SRAM
XU130 n45 n52 wordline[21] NOR2xp67_ASAP7_75t_SRAM
XU131 n45 n54 wordline[61] NOR2xp67_ASAP7_75t_SRAM
XU132 n45 n57 wordline[29] NOR2xp67_ASAP7_75t_SRAM
XU133 n45 n53 wordline[13] NOR2xp67_ASAP7_75t_SRAM
XU134 n45 n56 wordline[37] NOR2xp67_ASAP7_75t_SRAM
XU135 n58 n53 wordline[11] NOR2xp67_ASAP7_75t_SRAM
XU136 n58 n52 wordline[19] NOR2xp67_ASAP7_75t_SRAM
XU137 n58 n57 wordline[27] NOR2xp67_ASAP7_75t_SRAM
XU138 n58 n56 wordline[35] NOR2xp67_ASAP7_75t_SRAM
XU139 n58 n51 wordline[51] NOR2xp67_ASAP7_75t_SRAM
XU140 n58 n54 wordline[59] NOR2xp67_ASAP7_75t_SRAM
XU141 n47 n57 wordline[24] NOR2xp67_ASAP7_75t_SRAM
XU142 n47 n53 wordline[8] NOR2xp67_ASAP7_75t_SRAM
XU143 n47 n56 wordline[32] NOR2xp67_ASAP7_75t_SRAM
XU144 n47 n52 wordline[16] NOR2xp67_ASAP7_75t_SRAM
XU145 n47 n54 wordline[56] NOR2xp67_ASAP7_75t_SRAM
XU146 n47 n55 wordline[40] NOR2xp67_ASAP7_75t_SRAM
XU147 n47 n61 wordline[0] NOR2xp67_ASAP7_75t_SRAM
XU148 n47 n51 wordline[48] NOR2xp67_ASAP7_75t_SRAM
XU149 n59 n52 wordline[17] NOR2xp67_ASAP7_75t_SRAM
XU150 n59 n56 wordline[33] NOR2xp67_ASAP7_75t_SRAM
XU151 n59 n51 wordline[49] NOR2xp67_ASAP7_75t_SRAM
XU152 n60 n51 wordline[50] NOR2xp67_ASAP7_75t_SRAM
XU153 n59 n57 wordline[25] NOR2xp67_ASAP7_75t_SRAM
XU154 n60 n54 wordline[58] NOR2xp67_ASAP7_75t_SRAM
XU155 n60 n55 wordline[42] NOR2xp67_ASAP7_75t_SRAM
XU156 n60 n52 wordline[18] NOR2xp67_ASAP7_75t_SRAM
XU157 n60 n53 wordline[10] NOR2xp67_ASAP7_75t_SRAM
XU158 n59 n53 wordline[9] NOR2xp67_ASAP7_75t_SRAM
XU159 n59 n54 wordline[57] NOR2xp67_ASAP7_75t_SRAM
XU160 n59 n55 wordline[41] NOR2xp67_ASAP7_75t_SRAM
XU161 n60 n57 wordline[26] NOR2xp67_ASAP7_75t_SRAM
XU162 n61 n58 wordline[3] NOR2xp67_ASAP7_75t_SRAM
XU163 n61 n59 wordline[1] NOR2xp67_ASAP7_75t_SRAM
XU164 n61 n60 wordline[2] NOR2xp67_ASAP7_75t_SRAM
XU165 n42 n54 wordline[63] NOR2xp67_ASAP7_75t_SRAM
XU166 n43 n51 wordline[54] NOR2xp67_ASAP7_75t_SRAM
XU167 n58 n55 wordline[43] NOR2xp67_ASAP7_75t_SRAM
XU168 n60 n56 wordline[34] NOR2xp67_ASAP7_75t_SRAM
XU169 in_addr[5] n35 INVx5_ASAP7_75t_SRAM
XU170 in_addr[5] n36 INVx5_ASAP7_75t_SRAM
XU171 in_addr[5] n41 INVx5_ASAP7_75t_SRAM
XU172 in_addr[1] n37 INVx5_ASAP7_75t_SRAM
XU173 in_addr[1] n38 INVx5_ASAP7_75t_SRAM
XU174 in_addr[1] n48 INVx5_ASAP7_75t_SRAM
XU175 n35 n33 n39 n61 NAND3xp33_ASAP7_75t_SRAM
XU176 in_addr[1] clk in_addr[2] n49 n43 NAND4xp25_ASAP7_75t_SRAM
XU177 in_addr[0] clk in_addr[2] n48 n45 NAND4xp25_ASAP7_75t_SRAM
XU178 clk n28 n24 in_addr[2] n44 NAND4xp25_ASAP7_75t_SRAM
XU179 in_addr[0] in_addr[1] clk in_addr[2] n42 NAND4xp25_ASAP7_75t_SRAM
XU180 in_addr[4] in_addr[5] n25 n51 NAND3xp33_ASAP7_75t_SRAM
XU181 in_addr[5] in_addr[3] n26 n55 NAND3xp33_ASAP7_75t_SRAM
XU182 in_addr[5] n34 n29 n56 NAND3xp33_ASAP7_75t_SRAM
XU183 in_addr[5] in_addr[4] in_addr[3] n54 NAND3xp33_ASAP7_75t_SRAM
XU184 in_addr[4] n30 n27 n52 NAND3xp33_ASAP7_75t_SRAM
XU185 in_addr[3] n36 n40 n53 NAND3xp33_ASAP7_75t_SRAM
XU186 in_addr[4] in_addr[3] n41 n57 NAND3xp33_ASAP7_75t_SRAM
XU187 n46 in_addr[2] n50 NOR2xp33_ASAP7_75t_SRAM
XU188 in_addr[0] in_addr[1] n50 n58 NAND3xp33_ASAP7_75t_SRAM
XU189 n31 n37 n50 n47 NAND3xp33_ASAP7_75t_SRAM
XU190 in_addr[0] n50 n38 n59 NAND3xp33_ASAP7_75t_SRAM
XU191 in_addr[1] n50 n32 n60 NAND3xp33_ASAP7_75t_SRAM
.ENDS


